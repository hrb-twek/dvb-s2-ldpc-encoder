`timescale 1ns / 1ps
module enc_tbl_64800(
    clk,
    addr,
    dout
);
input wire clk;
input wire [13-1:0]addr;
output reg [20-1:0]dout;
always@(posedge clk) begin
    case(addr)
        default:  dout <= 0;
        // Q=135, BaseAddr=0
        'd0000: dout <= { 2'd1, 8'd116, 10'd174 }; 
        'd0001: dout <= { 2'd1, 8'd053, 10'd267 }; 
        'd0002: dout <= { 2'd1, 8'd060, 10'd008 }; 
        'd0003: dout <= { 2'd1, 8'd104, 10'd213 }; 
        'd0004: dout <= { 2'd1, 8'd058, 10'd134 }; 
        'd0005: dout <= { 2'd1, 8'd015, 10'd137 }; 
        'd0006: dout <= { 2'd1, 8'd016, 10'd046 }; 
        'd0007: dout <= { 2'd1, 8'd000, 10'd004 }; 
        'd0008: dout <= { 2'd1, 8'd029, 10'd311 }; 
        'd0009: dout <= { 2'd1, 8'd089, 10'd154 }; 
        'd0010: dout <= { 2'd1, 8'd042, 10'd176 }; 
        'd0011: dout <= { 2'd2, 8'd108, 10'd348 }; 
        'd0012: dout <= { 2'd1, 8'd084, 10'd121 }; 
        'd0013: dout <= { 2'd1, 8'd088, 10'd184 }; 
        'd0014: dout <= { 2'd1, 8'd004, 10'd123 }; 
        'd0015: dout <= { 2'd1, 8'd103, 10'd127 }; 
        'd0016: dout <= { 2'd1, 8'd133, 10'd056 }; 
        'd0017: dout <= { 2'd1, 8'd022, 10'd185 }; 
        'd0018: dout <= { 2'd1, 8'd062, 10'd315 }; 
        'd0019: dout <= { 2'd1, 8'd118, 10'd124 }; 
        'd0020: dout <= { 2'd1, 8'd091, 10'd258 }; 
        'd0021: dout <= { 2'd1, 8'd117, 10'd155 }; 
        'd0022: dout <= { 2'd1, 8'd034, 10'd274 }; 
        'd0023: dout <= { 2'd2, 8'd037, 10'd153 }; 
        'd0024: dout <= { 2'd1, 8'd119, 10'd013 }; 
        'd0025: dout <= { 2'd1, 8'd134, 10'd296 }; 
        'd0026: dout <= { 2'd1, 8'd074, 10'd138 }; 
        'd0027: dout <= { 2'd1, 8'd029, 10'd107 }; 
        'd0028: dout <= { 2'd1, 8'd099, 10'd103 }; 
        'd0029: dout <= { 2'd1, 8'd044, 10'd085 }; 
        'd0030: dout <= { 2'd1, 8'd011, 10'd097 }; 
        'd0031: dout <= { 2'd1, 8'd071, 10'd213 }; 
        'd0032: dout <= { 2'd1, 8'd059, 10'd286 }; 
        'd0033: dout <= { 2'd1, 8'd088, 10'd165 }; 
        'd0034: dout <= { 2'd1, 8'd015, 10'd224 }; 
        'd0035: dout <= { 2'd2, 8'd055, 10'd230 }; 
        'd0036: dout <= { 2'd1, 8'd114, 10'd164 }; 
        'd0037: dout <= { 2'd1, 8'd064, 10'd300 }; 
        'd0038: dout <= { 2'd1, 8'd100, 10'd167 }; 
        'd0039: dout <= { 2'd1, 8'd122, 10'd166 }; 
        'd0040: dout <= { 2'd1, 8'd059, 10'd045 }; 
        'd0041: dout <= { 2'd1, 8'd131, 10'd067 }; 
        'd0042: dout <= { 2'd1, 8'd038, 10'd296 }; 
        'd0043: dout <= { 2'd1, 8'd132, 10'd176 }; 
        'd0044: dout <= { 2'd1, 8'd027, 10'd066 }; 
        'd0045: dout <= { 2'd1, 8'd083, 10'd115 }; 
        'd0046: dout <= { 2'd1, 8'd114, 10'd124 }; 
        'd0047: dout <= { 2'd2, 8'd094, 10'd229 }; 
        'd0048: dout <= { 2'd1, 8'd072, 10'd059 }; 
        'd0049: dout <= { 2'd1, 8'd036, 10'd299 }; 
        'd0050: dout <= { 2'd1, 8'd050, 10'd100 }; 
        'd0051: dout <= { 2'd1, 8'd086, 10'd144 }; 
        'd0052: dout <= { 2'd1, 8'd052, 10'd310 }; 
        'd0053: dout <= { 2'd1, 8'd027, 10'd213 }; 
        'd0054: dout <= { 2'd1, 8'd074, 10'd098 }; 
        'd0055: dout <= { 2'd1, 8'd126, 10'd242 }; 
        'd0056: dout <= { 2'd1, 8'd109, 10'd182 }; 
        'd0057: dout <= { 2'd1, 8'd005, 10'd201 }; 
        'd0058: dout <= { 2'd1, 8'd080, 10'd340 }; 
        'd0059: dout <= { 2'd2, 8'd031, 10'd074 }; 
        'd0060: dout <= { 2'd1, 8'd040, 10'd300 }; 
        'd0061: dout <= { 2'd1, 8'd083, 10'd329 }; 
        'd0062: dout <= { 2'd1, 8'd006, 10'd103 }; 
        'd0063: dout <= { 2'd1, 8'd025, 10'd166 }; 
        'd0064: dout <= { 2'd1, 8'd031, 10'd242 }; 
        'd0065: dout <= { 2'd1, 8'd045, 10'd136 }; 
        'd0066: dout <= { 2'd1, 8'd104, 10'd295 }; 
        'd0067: dout <= { 2'd1, 8'd006, 10'd189 }; 
        'd0068: dout <= { 2'd1, 8'd077, 10'd092 }; 
        'd0069: dout <= { 2'd1, 8'd131, 10'd072 }; 
        'd0070: dout <= { 2'd1, 8'd073, 10'd290 }; 
        'd0071: dout <= { 2'd2, 8'd128, 10'd257 }; 
        'd0072: dout <= { 2'd1, 8'd113, 10'd112 }; 
        'd0073: dout <= { 2'd1, 8'd108, 10'd335 }; 
        'd0074: dout <= { 2'd1, 8'd046, 10'd037 }; 
        'd0075: dout <= { 2'd1, 8'd024, 10'd333 }; 
        'd0076: dout <= { 2'd1, 8'd080, 10'd338 }; 
        'd0077: dout <= { 2'd1, 8'd030, 10'd312 }; 
        'd0078: dout <= { 2'd1, 8'd111, 10'd143 }; 
        'd0079: dout <= { 2'd1, 8'd002, 10'd014 }; 
        'd0080: dout <= { 2'd1, 8'd036, 10'd171 }; 
        'd0081: dout <= { 2'd1, 8'd065, 10'd117 }; 
        'd0082: dout <= { 2'd1, 8'd057, 10'd065 }; 
        'd0083: dout <= { 2'd2, 8'd048, 10'd076 }; 
        'd0084: dout <= { 2'd1, 8'd073, 10'd077 }; 
        'd0085: dout <= { 2'd1, 8'd016, 10'd328 }; 
        'd0086: dout <= { 2'd1, 8'd101, 10'd026 }; 
        'd0087: dout <= { 2'd1, 8'd130, 10'd010 }; 
        'd0088: dout <= { 2'd1, 8'd051, 10'd278 }; 
        'd0089: dout <= { 2'd1, 8'd124, 10'd238 }; 
        'd0090: dout <= { 2'd1, 8'd047, 10'd102 }; 
        'd0091: dout <= { 2'd1, 8'd133, 10'd050 }; 
        'd0092: dout <= { 2'd1, 8'd087, 10'd243 }; 
        'd0093: dout <= { 2'd1, 8'd028, 10'd298 }; 
        'd0094: dout <= { 2'd1, 8'd098, 10'd344 }; 
        'd0095: dout <= { 2'd2, 8'd060, 10'd088 }; 
        'd0096: dout <= { 2'd1, 8'd090, 10'd049 }; 
        'd0097: dout <= { 2'd1, 8'd034, 10'd160 }; 
        'd0098: dout <= { 2'd1, 8'd070, 10'd208 }; 
        'd0099: dout <= { 2'd1, 8'd017, 10'd324 }; 
        'd0100: dout <= { 2'd1, 8'd085, 10'd006 }; 
        'd0101: dout <= { 2'd1, 8'd067, 10'd048 }; 
        'd0102: dout <= { 2'd1, 8'd045, 10'd155 }; 
        'd0103: dout <= { 2'd1, 8'd024, 10'd214 }; 
        'd0104: dout <= { 2'd1, 8'd012, 10'd223 }; 
        'd0105: dout <= { 2'd1, 8'd086, 10'd190 }; 
        'd0106: dout <= { 2'd1, 8'd019, 10'd309 }; 
        'd0107: dout <= { 2'd2, 8'd052, 10'd084 }; 
        'd0108: dout <= { 2'd1, 8'd132, 10'd162 }; 
        'd0109: dout <= { 2'd1, 8'd069, 10'd042 }; 
        'd0110: dout <= { 2'd1, 8'd075, 10'd201 }; 
        'd0111: dout <= { 2'd1, 8'd018, 10'd206 }; 
        'd0112: dout <= { 2'd1, 8'd037, 10'd253 }; 
        'd0113: dout <= { 2'd1, 8'd057, 10'd281 }; 
        'd0114: dout <= { 2'd1, 8'd115, 10'd080 }; 
        'd0115: dout <= { 2'd1, 8'd113, 10'd051 }; 
        'd0116: dout <= { 2'd1, 8'd044, 10'd028 }; 
        'd0117: dout <= { 2'd1, 8'd010, 10'd312 }; 
        'd0118: dout <= { 2'd1, 8'd039, 10'd033 }; 
        'd0119: dout <= { 2'd2, 8'd099, 10'd264 }; 
        'd0120: dout <= { 2'd1, 8'd010, 10'd063 }; 
        'd0121: dout <= { 2'd1, 8'd111, 10'd008 }; 
        'd0122: dout <= { 2'd1, 8'd007, 10'd101 }; 
        'd0123: dout <= { 2'd1, 8'd035, 10'd229 }; 
        'd0124: dout <= { 2'd1, 8'd023, 10'd192 }; 
        'd0125: dout <= { 2'd1, 8'd118, 10'd093 }; 
        'd0126: dout <= { 2'd1, 8'd121, 10'd123 }; 
        'd0127: dout <= { 2'd1, 8'd106, 10'd253 }; 
        'd0128: dout <= { 2'd1, 8'd103, 10'd235 }; 
        'd0129: dout <= { 2'd1, 8'd100, 10'd024 }; 
        'd0130: dout <= { 2'd1, 8'd107, 10'd064 }; 
        'd0131: dout <= { 2'd2, 8'd075, 10'd290 }; 
        'd0132: dout <= { 2'd1, 8'd079, 10'd140 }; 
        'd0133: dout <= { 2'd1, 8'd048, 10'd126 }; 
        'd0134: dout <= { 2'd1, 8'd065, 10'd319 }; 
        'd0135: dout <= { 2'd1, 8'd061, 10'd031 }; 
        'd0136: dout <= { 2'd1, 8'd068, 10'd035 }; 
        'd0137: dout <= { 2'd1, 8'd020, 10'd326 }; 
        'd0138: dout <= { 2'd1, 8'd014, 10'd144 }; 
        'd0139: dout <= { 2'd1, 8'd081, 10'd218 }; 
        'd0140: dout <= { 2'd1, 8'd004, 10'd355 }; 
        'd0141: dout <= { 2'd1, 8'd054, 10'd112 }; 
        'd0142: dout <= { 2'd1, 8'd033, 10'd180 }; 
        'd0143: dout <= { 2'd2, 8'd049, 10'd143 }; 
        'd0144: dout <= { 2'd1, 8'd089, 10'd123 }; 
        'd0145: dout <= { 2'd1, 8'd011, 10'd062 }; 
        'd0146: dout <= { 2'd1, 8'd077, 10'd219 }; 
        'd0147: dout <= { 2'd1, 8'd076, 10'd344 }; 
        'd0148: dout <= { 2'd1, 8'd094, 10'd238 }; 
        'd0149: dout <= { 2'd1, 8'd019, 10'd195 }; 
        'd0150: dout <= { 2'd1, 8'd090, 10'd069 }; 
        'd0151: dout <= { 2'd1, 8'd067, 10'd135 }; 
        'd0152: dout <= { 2'd1, 8'd017, 10'd092 }; 
        'd0153: dout <= { 2'd1, 8'd046, 10'd202 }; 
        'd0154: dout <= { 2'd1, 8'd096, 10'd262 }; 
        'd0155: dout <= { 2'd2, 8'd007, 10'd311 }; 
        'd0156: dout <= { 2'd1, 8'd117, 10'd115 }; 
        'd0157: dout <= { 2'd1, 8'd066, 10'd043 }; 
        'd0158: dout <= { 2'd1, 8'd049, 10'd344 }; 
        'd0159: dout <= { 2'd1, 8'd128, 10'd197 }; 
        'd0160: dout <= { 2'd1, 8'd041, 10'd173 }; 
        'd0161: dout <= { 2'd1, 8'd102, 10'd053 }; 
        'd0162: dout <= { 2'd1, 8'd064, 10'd066 }; 
        'd0163: dout <= { 2'd1, 8'd051, 10'd023 }; 
        'd0164: dout <= { 2'd1, 8'd025, 10'd277 }; 
        'd0165: dout <= { 2'd1, 8'd003, 10'd332 }; 
        'd0166: dout <= { 2'd1, 8'd053, 10'd262 }; 
        'd0167: dout <= { 2'd2, 8'd041, 10'd100 }; 
        'd0168: dout <= { 2'd1, 8'd063, 10'd317 }; 
        'd0169: dout <= { 2'd1, 8'd013, 10'd237 }; 
        'd0170: dout <= { 2'd1, 8'd107, 10'd305 }; 
        'd0171: dout <= { 2'd1, 8'd028, 10'd287 }; 
        'd0172: dout <= { 2'd1, 8'd110, 10'd196 }; 
        'd0173: dout <= { 2'd1, 8'd002, 10'd020 }; 
        'd0174: dout <= { 2'd1, 8'd125, 10'd201 }; 
        'd0175: dout <= { 2'd1, 8'd129, 10'd347 }; 
        'd0176: dout <= { 2'd1, 8'd119, 10'd010 }; 
        'd0177: dout <= { 2'd1, 8'd097, 10'd154 }; 
        'd0178: dout <= { 2'd1, 8'd021, 10'd203 }; 
        'd0179: dout <= { 2'd2, 8'd078, 10'd285 }; 
        'd0180: dout <= { 2'd1, 8'd012, 10'd164 }; 
        'd0181: dout <= { 2'd1, 8'd096, 10'd179 }; 
        'd0182: dout <= { 2'd2, 8'd062, 10'd061 }; 
        'd0183: dout <= { 2'd1, 8'd042, 10'd143 }; 
        'd0184: dout <= { 2'd1, 8'd123, 10'd073 }; 
        'd0185: dout <= { 2'd2, 8'd127, 10'd205 }; 
        'd0186: dout <= { 2'd1, 8'd026, 10'd259 }; 
        'd0187: dout <= { 2'd1, 8'd009, 10'd047 }; 
        'd0188: dout <= { 2'd2, 8'd081, 10'd248 }; 
        'd0189: dout <= { 2'd1, 8'd082, 10'd220 }; 
        'd0190: dout <= { 2'd1, 8'd095, 10'd228 }; 
        'd0191: dout <= { 2'd2, 8'd093, 10'd218 }; 
        'd0192: dout <= { 2'd1, 8'd098, 10'd068 }; 
        'd0193: dout <= { 2'd1, 8'd047, 10'd359 }; 
        'd0194: dout <= { 2'd2, 8'd039, 10'd106 }; 
        'd0195: dout <= { 2'd1, 8'd126, 10'd281 }; 
        'd0196: dout <= { 2'd1, 8'd115, 10'd030 }; 
        'd0197: dout <= { 2'd2, 8'd003, 10'd325 }; 
        'd0198: dout <= { 2'd1, 8'd043, 10'd063 }; 
        'd0199: dout <= { 2'd1, 8'd097, 10'd245 }; 
        'd0200: dout <= { 2'd2, 8'd120, 10'd254 }; 
        'd0201: dout <= { 2'd1, 8'd125, 10'd166 }; 
        'd0202: dout <= { 2'd1, 8'd056, 10'd213 }; 
        'd0203: dout <= { 2'd2, 8'd055, 10'd177 }; 
        'd0204: dout <= { 2'd1, 8'd054, 10'd151 }; 
        'd0205: dout <= { 2'd1, 8'd112, 10'd029 }; 
        'd0206: dout <= { 2'd2, 8'd021, 10'd179 }; 
        'd0207: dout <= { 2'd1, 8'd008, 10'd286 }; 
        'd0208: dout <= { 2'd1, 8'd087, 10'd060 }; 
        'd0209: dout <= { 2'd2, 8'd032, 10'd229 }; 
        'd0210: dout <= { 2'd1, 8'd033, 10'd263 }; 
        'd0211: dout <= { 2'd1, 8'd005, 10'd325 }; 
        'd0212: dout <= { 2'd2, 8'd129, 10'd158 }; 
        'd0213: dout <= { 2'd1, 8'd071, 10'd052 }; 
        'd0214: dout <= { 2'd1, 8'd121, 10'd337 }; 
        'd0215: dout <= { 2'd2, 8'd078, 10'd111 }; 
        'd0216: dout <= { 2'd1, 8'd105, 10'd040 }; 
        'd0217: dout <= { 2'd1, 8'd000, 10'd069 }; 
        'd0218: dout <= { 2'd2, 8'd038, 10'd162 }; 
        'd0219: dout <= { 2'd1, 8'd001, 10'd267 }; 
        'd0220: dout <= { 2'd1, 8'd109, 10'd243 }; 
        'd0221: dout <= { 2'd2, 8'd091, 10'd087 }; 
        'd0222: dout <= { 2'd1, 8'd014, 10'd054 }; 
        'd0223: dout <= { 2'd1, 8'd092, 10'd294 }; 
        'd0224: dout <= { 2'd2, 8'd106, 10'd249 }; 
        'd0225: dout <= { 2'd1, 8'd030, 10'd125 }; 
        'd0226: dout <= { 2'd1, 8'd127, 10'd221 }; 
        'd0227: dout <= { 2'd2, 8'd020, 10'd096 }; 
        'd0228: dout <= { 2'd1, 8'd101, 10'd082 }; 
        'd0229: dout <= { 2'd1, 8'd084, 10'd175 }; 
        'd0230: dout <= { 2'd2, 8'd050, 10'd166 }; 
        'd0231: dout <= { 2'd1, 8'd116, 10'd255 }; 
        'd0232: dout <= { 2'd1, 8'd082, 10'd073 }; 
        'd0233: dout <= { 2'd2, 8'd085, 10'd329 }; 
        'd0234: dout <= { 2'd1, 8'd130, 10'd103 }; 
        'd0235: dout <= { 2'd1, 8'd066, 10'd350 }; 
        'd0236: dout <= { 2'd2, 8'd040, 10'd065 }; 
        'd0237: dout <= { 2'd1, 8'd072, 10'd111 }; 
        'd0238: dout <= { 2'd1, 8'd122, 10'd336 }; 
        'd0239: dout <= { 2'd2, 8'd026, 10'd181 }; 
        'd0240: dout <= { 2'd1, 8'd008, 10'd226 }; 
        'd0241: dout <= { 2'd1, 8'd022, 10'd273 }; 
        'd0242: dout <= { 2'd2, 8'd069, 10'd006 }; 
        'd0243: dout <= { 2'd1, 8'd023, 10'd056 }; 
        'd0244: dout <= { 2'd1, 8'd134, 10'd098 }; 
        'd0245: dout <= { 2'd2, 8'd032, 10'd180 }; 
        'd0246: dout <= { 2'd1, 8'd043, 10'd003 }; 
        'd0247: dout <= { 2'd1, 8'd056, 10'd200 }; 
        'd0248: dout <= { 2'd2, 8'd092, 10'd034 }; 
        'd0249: dout <= { 2'd1, 8'd068, 10'd089 }; 
        'd0250: dout <= { 2'd1, 8'd058, 10'd232 }; 
        'd0251: dout <= { 2'd2, 8'd070, 10'd160 }; 
        'd0252: dout <= { 2'd1, 8'd079, 10'd008 }; 
        'd0253: dout <= { 2'd1, 8'd076, 10'd133 }; 
        'd0254: dout <= { 2'd2, 8'd061, 10'd016 }; 
        'd0255: dout <= { 2'd1, 8'd018, 10'd126 }; 
        'd0256: dout <= { 2'd1, 8'd105, 10'd286 }; 
        'd0257: dout <= { 2'd2, 8'd035, 10'd069 }; 
        'd0258: dout <= { 2'd1, 8'd063, 10'd128 }; 
        'd0259: dout <= { 2'd1, 8'd095, 10'd181 }; 
        'd0260: dout <= { 2'd2, 8'd009, 10'd219 }; 
        'd0261: dout <= { 2'd1, 8'd093, 10'd341 }; 
        'd0262: dout <= { 2'd1, 8'd124, 10'd229 }; 
        'd0263: dout <= { 2'd2, 8'd013, 10'd243 }; 
        'd0264: dout <= { 2'd1, 8'd123, 10'd150 }; 
        'd0265: dout <= { 2'd1, 8'd112, 10'd273 }; 
        'd0266: dout <= { 2'd2, 8'd120, 10'd135 }; 
        'd0267: dout <= { 2'd1, 8'd110, 10'd345 }; 
        'd0268: dout <= { 2'd1, 8'd102, 10'd152 }; 
        'd0269: dout <= { 2'd3, 8'd001, 10'd243 }; 
        // Q=120, BaseAddr=270
        'd0270: dout <= { 2'd1, 8'd103, 10'd290 }; 
        'd0271: dout <= { 2'd1, 8'd047, 10'd174 }; 
        'd0272: dout <= { 2'd1, 8'd053, 10'd267 }; 
        'd0273: dout <= { 2'd1, 8'd092, 10'd008 }; 
        'd0274: dout <= { 2'd1, 8'd051, 10'd213 }; 
        'd0275: dout <= { 2'd1, 8'd013, 10'd134 }; 
        'd0276: dout <= { 2'd1, 8'd014, 10'd137 }; 
        'd0277: dout <= { 2'd1, 8'd000, 10'd046 }; 
        'd0278: dout <= { 2'd1, 8'd026, 10'd004 }; 
        'd0279: dout <= { 2'd1, 8'd079, 10'd311 }; 
        'd0280: dout <= { 2'd1, 8'd038, 10'd154 }; 
        'd0281: dout <= { 2'd2, 8'd000, 10'd176 }; 
        'd0282: dout <= { 2'd1, 8'd116, 10'd096 }; 
        'd0283: dout <= { 2'd1, 8'd074, 10'd121 }; 
        'd0284: dout <= { 2'd1, 8'd078, 10'd184 }; 
        'd0285: dout <= { 2'd1, 8'd003, 10'd123 }; 
        'd0286: dout <= { 2'd1, 8'd093, 10'd127 }; 
        'd0287: dout <= { 2'd1, 8'd118, 10'd056 }; 
        'd0288: dout <= { 2'd1, 8'd022, 10'd185 }; 
        'd0289: dout <= { 2'd1, 8'd056, 10'd315 }; 
        'd0290: dout <= { 2'd1, 8'd105, 10'd124 }; 
        'd0291: dout <= { 2'd1, 8'd081, 10'd258 }; 
        'd0292: dout <= { 2'd1, 8'd104, 10'd155 }; 
        'd0293: dout <= { 2'd2, 8'd030, 10'd274 }; 
        'd0294: dout <= { 2'd1, 8'd049, 10'd145 }; 
        'd0295: dout <= { 2'd1, 8'd105, 10'd013 }; 
        'd0296: dout <= { 2'd1, 8'd119, 10'd296 }; 
        'd0297: dout <= { 2'd1, 8'd064, 10'd138 }; 
        'd0298: dout <= { 2'd1, 8'd027, 10'd107 }; 
        'd0299: dout <= { 2'd1, 8'd089, 10'd103 }; 
        'd0300: dout <= { 2'd1, 8'd041, 10'd085 }; 
        'd0301: dout <= { 2'd1, 8'd010, 10'd097 }; 
        'd0302: dout <= { 2'd1, 8'd062, 10'd213 }; 
        'd0303: dout <= { 2'd1, 8'd052, 10'd286 }; 
        'd0304: dout <= { 2'd1, 8'd078, 10'd165 }; 
        'd0305: dout <= { 2'd2, 8'd014, 10'd224 }; 
        'd0306: dout <= { 2'd1, 8'd075, 10'd243 }; 
        'd0307: dout <= { 2'd1, 8'd100, 10'd164 }; 
        'd0308: dout <= { 2'd1, 8'd056, 10'd300 }; 
        'd0309: dout <= { 2'd1, 8'd089, 10'd167 }; 
        'd0310: dout <= { 2'd1, 8'd109, 10'd166 }; 
        'd0311: dout <= { 2'd1, 8'd057, 10'd045 }; 
        'd0312: dout <= { 2'd1, 8'd117, 10'd067 }; 
        'd0313: dout <= { 2'd1, 8'd034, 10'd296 }; 
        'd0314: dout <= { 2'd1, 8'd117, 10'd176 }; 
        'd0315: dout <= { 2'd1, 8'd023, 10'd066 }; 
        'd0316: dout <= { 2'd1, 8'd073, 10'd115 }; 
        'd0317: dout <= { 2'd2, 8'd100, 10'd124 }; 
        'd0318: dout <= { 2'd1, 8'd072, 10'd082 }; 
        'd0319: dout <= { 2'd1, 8'd063, 10'd059 }; 
        'd0320: dout <= { 2'd1, 8'd031, 10'd299 }; 
        'd0321: dout <= { 2'd1, 8'd043, 10'd100 }; 
        'd0322: dout <= { 2'd1, 8'd080, 10'd144 }; 
        'd0323: dout <= { 2'd1, 8'd053, 10'd310 }; 
        'd0324: dout <= { 2'd1, 8'd028, 10'd213 }; 
        'd0325: dout <= { 2'd1, 8'd067, 10'd098 }; 
        'd0326: dout <= { 2'd1, 8'd112, 10'd242 }; 
        'd0327: dout <= { 2'd1, 8'd096, 10'd182 }; 
        'd0328: dout <= { 2'd1, 8'd005, 10'd201 }; 
        'd0329: dout <= { 2'd2, 8'd070, 10'd340 }; 
        'd0330: dout <= { 2'd1, 8'd021, 10'd339 }; 
        'd0331: dout <= { 2'd1, 8'd035, 10'd300 }; 
        'd0332: dout <= { 2'd1, 8'd076, 10'd329 }; 
        'd0333: dout <= { 2'd1, 8'd006, 10'd103 }; 
        'd0334: dout <= { 2'd1, 8'd026, 10'd166 }; 
        'd0335: dout <= { 2'd1, 8'd032, 10'd242 }; 
        'd0336: dout <= { 2'd1, 8'd045, 10'd136 }; 
        'd0337: dout <= { 2'd1, 8'd095, 10'd295 }; 
        'd0338: dout <= { 2'd1, 8'd006, 10'd189 }; 
        'd0339: dout <= { 2'd1, 8'd066, 10'd092 }; 
        'd0340: dout <= { 2'd1, 8'd116, 10'd072 }; 
        'd0341: dout <= { 2'd2, 8'd063, 10'd290 }; 
        'd0342: dout <= { 2'd1, 8'd085, 10'd159 }; 
        'd0343: dout <= { 2'd1, 8'd102, 10'd130 }; 
        'd0344: dout <= { 2'd1, 8'd096, 10'd112 }; 
        'd0345: dout <= { 2'd1, 8'd038, 10'd335 }; 
        'd0346: dout <= { 2'd1, 8'd025, 10'd037 }; 
        'd0347: dout <= { 2'd1, 8'd074, 10'd333 }; 
        'd0348: dout <= { 2'd1, 8'd030, 10'd338 }; 
        'd0349: dout <= { 2'd1, 8'd100, 10'd312 }; 
        'd0350: dout <= { 2'd1, 8'd002, 10'd143 }; 
        'd0351: dout <= { 2'd1, 8'd032, 10'd014 }; 
        'd0352: dout <= { 2'd1, 8'd057, 10'd171 }; 
        'd0353: dout <= { 2'd2, 8'd098, 10'd117 }; 
        'd0354: dout <= { 2'd1, 8'd018, 10'd261 }; 
        'd0355: dout <= { 2'd1, 8'd022, 10'd161 }; 
        'd0356: dout <= { 2'd1, 8'd061, 10'd077 }; 
        'd0357: dout <= { 2'd1, 8'd015, 10'd328 }; 
        'd0358: dout <= { 2'd1, 8'd091, 10'd026 }; 
        'd0359: dout <= { 2'd1, 8'd116, 10'd010 }; 
        'd0360: dout <= { 2'd1, 8'd049, 10'd278 }; 
        'd0361: dout <= { 2'd1, 8'd110, 10'd238 }; 
        'd0362: dout <= { 2'd1, 8'd042, 10'd102 }; 
        'd0363: dout <= { 2'd1, 8'd118, 10'd050 }; 
        'd0364: dout <= { 2'd1, 8'd076, 10'd243 }; 
        'd0365: dout <= { 2'd2, 8'd027, 10'd298 }; 
        'd0366: dout <= { 2'd1, 8'd104, 10'd095 }; 
        'd0367: dout <= { 2'd1, 8'd026, 10'd254 }; 
        'd0368: dout <= { 2'd1, 8'd118, 10'd162 }; 
        'd0369: dout <= { 2'd1, 8'd060, 10'd042 }; 
        'd0370: dout <= { 2'd1, 8'd068, 10'd201 }; 
        'd0371: dout <= { 2'd1, 8'd018, 10'd206 }; 
        'd0372: dout <= { 2'd1, 8'd037, 10'd253 }; 
        'd0373: dout <= { 2'd1, 8'd055, 10'd281 }; 
        'd0374: dout <= { 2'd1, 8'd099, 10'd080 }; 
        'd0375: dout <= { 2'd1, 8'd095, 10'd051 }; 
        'd0376: dout <= { 2'd1, 8'd037, 10'd028 }; 
        'd0377: dout <= { 2'd2, 8'd011, 10'd312 }; 
        'd0378: dout <= { 2'd1, 8'd009, 10'd289 }; 
        'd0379: dout <= { 2'd1, 8'd086, 10'd192 }; 
        'd0380: dout <= { 2'd1, 8'd011, 10'd063 }; 
        'd0381: dout <= { 2'd1, 8'd098, 10'd008 }; 
        'd0382: dout <= { 2'd1, 8'd007, 10'd101 }; 
        'd0383: dout <= { 2'd1, 8'd038, 10'd229 }; 
        'd0384: dout <= { 2'd1, 8'd024, 10'd192 }; 
        'd0385: dout <= { 2'd1, 8'd105, 10'd093 }; 
        'd0386: dout <= { 2'd1, 8'd107, 10'd123 }; 
        'd0387: dout <= { 2'd1, 8'd091, 10'd253 }; 
        'd0388: dout <= { 2'd1, 8'd089, 10'd235 }; 
        'd0389: dout <= { 2'd2, 8'd086, 10'd024 }; 
        'd0390: dout <= { 2'd1, 8'd020, 10'd097 }; 
        'd0391: dout <= { 2'd1, 8'd094, 10'd127 }; 
        'd0392: dout <= { 2'd1, 8'd067, 10'd140 }; 
        'd0393: dout <= { 2'd1, 8'd040, 10'd126 }; 
        'd0394: dout <= { 2'd1, 8'd063, 10'd319 }; 
        'd0395: dout <= { 2'd1, 8'd058, 10'd031 }; 
        'd0396: dout <= { 2'd1, 8'd065, 10'd035 }; 
        'd0397: dout <= { 2'd1, 8'd019, 10'd326 }; 
        'd0398: dout <= { 2'd1, 8'd013, 10'd144 }; 
        'd0399: dout <= { 2'd1, 8'd069, 10'd218 }; 
        'd0400: dout <= { 2'd1, 8'd004, 10'd355 }; 
        'd0401: dout <= { 2'd2, 8'd046, 10'd112 }; 
        'd0402: dout <= { 2'd1, 8'd057, 10'd262 }; 
        'd0403: dout <= { 2'd1, 8'd045, 10'd011 }; 
        'd0404: dout <= { 2'd1, 8'd068, 10'd123 }; 
        'd0405: dout <= { 2'd1, 8'd013, 10'd062 }; 
        'd0406: dout <= { 2'd1, 8'd070, 10'd219 }; 
        'd0407: dout <= { 2'd1, 8'd066, 10'd344 }; 
        'd0408: dout <= { 2'd1, 8'd083, 10'd238 }; 
        'd0409: dout <= { 2'd1, 8'd021, 10'd195 }; 
        'd0410: dout <= { 2'd1, 8'd074, 10'd069 }; 
        'd0411: dout <= { 2'd1, 8'd055, 10'd135 }; 
        'd0412: dout <= { 2'd1, 8'd015, 10'd092 }; 
        'd0413: dout <= { 2'd2, 8'd039, 10'd202 }; 
        'd0414: dout <= { 2'd1, 8'd087, 10'd130 }; 
        'd0415: dout <= { 2'd1, 8'd107, 10'd103 }; 
        'd0416: dout <= { 2'd1, 8'd106, 10'd115 }; 
        'd0417: dout <= { 2'd1, 8'd055, 10'd043 }; 
        'd0418: dout <= { 2'd1, 8'd048, 10'd344 }; 
        'd0419: dout <= { 2'd1, 8'd115, 10'd197 }; 
        'd0420: dout <= { 2'd1, 8'd040, 10'd173 }; 
        'd0421: dout <= { 2'd1, 8'd087, 10'd053 }; 
        'd0422: dout <= { 2'd1, 8'd050, 10'd066 }; 
        'd0423: dout <= { 2'd1, 8'd043, 10'd023 }; 
        'd0424: dout <= { 2'd1, 8'd022, 10'd277 }; 
        'd0425: dout <= { 2'd2, 8'd003, 10'd332 }; 
        'd0426: dout <= { 2'd1, 8'd083, 10'd044 }; 
        'd0427: dout <= { 2'd1, 8'd029, 10'd187 }; 
        'd0428: dout <= { 2'd1, 8'd051, 10'd317 }; 
        'd0429: dout <= { 2'd1, 8'd017, 10'd237 }; 
        'd0430: dout <= { 2'd1, 8'd096, 10'd305 }; 
        'd0431: dout <= { 2'd1, 8'd031, 10'd287 }; 
        'd0432: dout <= { 2'd1, 8'd099, 10'd196 }; 
        'd0433: dout <= { 2'd1, 8'd004, 10'd020 }; 
        'd0434: dout <= { 2'd1, 8'd109, 10'd201 }; 
        'd0435: dout <= { 2'd1, 8'd114, 10'd347 }; 
        'd0436: dout <= { 2'd1, 8'd097, 10'd010 }; 
        'd0437: dout <= { 2'd2, 8'd083, 10'd154 }; 
        'd0438: dout <= { 2'd1, 8'd073, 10'd030 }; 
        'd0439: dout <= { 2'd1, 8'd070, 10'd325 }; 
        'd0440: dout <= { 2'd1, 8'd080, 10'd120 }; 
        'd0441: dout <= { 2'd1, 8'd039, 10'd252 }; 
        'd0442: dout <= { 2'd1, 8'd043, 10'd312 }; 
        'd0443: dout <= { 2'd1, 8'd020, 10'd063 }; 
        'd0444: dout <= { 2'd1, 8'd119, 10'd245 }; 
        'd0445: dout <= { 2'd1, 8'd039, 10'd254 }; 
        'd0446: dout <= { 2'd1, 8'd111, 10'd331 }; 
        'd0447: dout <= { 2'd1, 8'd092, 10'd168 }; 
        'd0448: dout <= { 2'd1, 8'd012, 10'd151 }; 
        'd0449: dout <= { 2'd2, 8'd090, 10'd166 }; 
        'd0450: dout <= { 2'd1, 8'd066, 10'd286 }; 
        'd0451: dout <= { 2'd1, 8'd052, 10'd060 }; 
        'd0452: dout <= { 2'd1, 8'd046, 10'd229 }; 
        'd0453: dout <= { 2'd1, 8'd110, 10'd107 }; 
        'd0454: dout <= { 2'd1, 8'd035, 10'd057 }; 
        'd0455: dout <= { 2'd1, 8'd060, 10'd358 }; 
        'd0456: dout <= { 2'd1, 8'd006, 10'd263 }; 
        'd0457: dout <= { 2'd1, 8'd069, 10'd325 }; 
        'd0458: dout <= { 2'd1, 8'd025, 10'd158 }; 
        'd0459: dout <= { 2'd1, 8'd061, 10'd129 }; 
        'd0460: dout <= { 2'd1, 8'd060, 10'd333 }; 
        'd0461: dout <= { 2'd2, 8'd035, 10'd139 }; 
        'd0462: dout <= { 2'd1, 8'd041, 10'd014 }; 
        'd0463: dout <= { 2'd1, 8'd012, 10'd311 }; 
        'd0464: dout <= { 2'd1, 8'd113, 10'd332 }; 
        'd0465: dout <= { 2'd1, 8'd030, 10'd145 }; 
        'd0466: dout <= { 2'd1, 8'd094, 10'd267 }; 
        'd0467: dout <= { 2'd1, 8'd002, 10'd243 }; 
        'd0468: dout <= { 2'd1, 8'd050, 10'd087 }; 
        'd0469: dout <= { 2'd1, 8'd011, 10'd108 }; 
        'd0470: dout <= { 2'd1, 8'd021, 10'd238 }; 
        'd0471: dout <= { 2'd1, 8'd051, 10'd244 }; 
        'd0472: dout <= { 2'd1, 8'd009, 10'd054 }; 
        'd0473: dout <= { 2'd2, 8'd103, 10'd294 }; 
        'd0474: dout <= { 2'd1, 8'd016, 10'd006 }; 
        'd0475: dout <= { 2'd1, 8'd062, 10'd058 }; 
        'd0476: dout <= { 2'd1, 8'd109, 10'd352 }; 
        'd0477: dout <= { 2'd1, 8'd023, 10'd073 }; 
        'd0478: dout <= { 2'd1, 8'd047, 10'd056 }; 
        'd0479: dout <= { 2'd1, 8'd111, 10'd098 }; 
        'd0480: dout <= { 2'd1, 8'd075, 10'd180 }; 
        'd0481: dout <= { 2'd1, 8'd005, 10'd086 }; 
        'd0482: dout <= { 2'd1, 8'd028, 10'd096 }; 
        'd0483: dout <= { 2'd1, 8'd058, 10'd216 }; 
        'd0484: dout <= { 2'd1, 8'd071, 10'd003 }; 
        'd0485: dout <= { 2'd2, 8'd085, 10'd200 }; 
        'd0486: dout <= { 2'd1, 8'd005, 10'd016 }; 
        'd0487: dout <= { 2'd1, 8'd042, 10'd088 }; 
        'd0488: dout <= { 2'd1, 8'd025, 10'd238 }; 
        'd0489: dout <= { 2'd1, 8'd050, 10'd101 }; 
        'd0490: dout <= { 2'd1, 8'd036, 10'd126 }; 
        'd0491: dout <= { 2'd1, 8'd084, 10'd286 }; 
        'd0492: dout <= { 2'd1, 8'd071, 10'd069 }; 
        'd0493: dout <= { 2'd1, 8'd073, 10'd110 }; 
        'd0494: dout <= { 2'd1, 8'd048, 10'd168 }; 
        'd0495: dout <= { 2'd1, 8'd040, 10'd048 }; 
        'd0496: dout <= { 2'd1, 8'd007, 10'd128 }; 
        'd0497: dout <= { 2'd2, 8'd044, 10'd181 }; 
        'd0498: dout <= { 2'd1, 8'd079, 10'd135 }; 
        'd0499: dout <= { 2'd1, 8'd032, 10'd315 }; 
        'd0500: dout <= { 2'd1, 8'd112, 10'd289 }; 
        'd0501: dout <= { 2'd1, 8'd010, 10'd177 }; 
        'd0502: dout <= { 2'd1, 8'd112, 10'd284 }; 
        'd0503: dout <= { 2'd1, 8'd086, 10'd061 }; 
        'd0504: dout <= { 2'd1, 8'd088, 10'd345 }; 
        'd0505: dout <= { 2'd1, 8'd106, 10'd152 }; 
        'd0506: dout <= { 2'd1, 8'd067, 10'd243 }; 
        'd0507: dout <= { 2'd1, 8'd087, 10'd217 }; 
        'd0508: dout <= { 2'd1, 8'd053, 10'd212 }; 
        'd0509: dout <= { 2'd2, 8'd088, 10'd058 }; 
        'd0510: dout <= { 2'd1, 8'd108, 10'd332 }; 
        'd0511: dout <= { 2'd1, 8'd029, 10'd235 }; 
        'd0512: dout <= { 2'd2, 8'd059, 10'd207 }; 
        'd0513: dout <= { 2'd1, 8'd008, 10'd145 }; 
        'd0514: dout <= { 2'd1, 8'd114, 10'd118 }; 
        'd0515: dout <= { 2'd2, 8'd113, 10'd324 }; 
        'd0516: dout <= { 2'd1, 8'd014, 10'd323 }; 
        'd0517: dout <= { 2'd1, 8'd008, 10'd133 }; 
        'd0518: dout <= { 2'd2, 8'd019, 10'd237 }; 
        'd0519: dout <= { 2'd1, 8'd004, 10'd345 }; 
        'd0520: dout <= { 2'd1, 8'd009, 10'd227 }; 
        'd0521: dout <= { 2'd2, 8'd065, 10'd228 }; 
        'd0522: dout <= { 2'd1, 8'd069, 10'd343 }; 
        'd0523: dout <= { 2'd1, 8'd082, 10'd050 }; 
        'd0524: dout <= { 2'd2, 8'd034, 10'd359 }; 
        'd0525: dout <= { 2'd1, 8'd037, 10'd116 }; 
        'd0526: dout <= { 2'd1, 8'd059, 10'd041 }; 
        'd0527: dout <= { 2'd2, 8'd094, 10'd338 }; 
        'd0528: dout <= { 2'd1, 8'd093, 10'd025 }; 
        'd0529: dout <= { 2'd1, 8'd078, 10'd028 }; 
        'd0530: dout <= { 2'd2, 8'd072, 10'd291 }; 
        'd0531: dout <= { 2'd1, 8'd002, 10'd284 }; 
        'd0532: dout <= { 2'd1, 8'd052, 10'd051 }; 
        'd0533: dout <= { 2'd2, 8'd080, 10'd239 }; 
        'd0534: dout <= { 2'd1, 8'd090, 10'd351 }; 
        'd0535: dout <= { 2'd1, 8'd061, 10'd284 }; 
        'd0536: dout <= { 2'd2, 8'd101, 10'd341 }; 
        'd0537: dout <= { 2'd1, 8'd065, 10'd122 }; 
        'd0538: dout <= { 2'd1, 8'd023, 10'd148 }; 
        'd0539: dout <= { 2'd2, 8'd054, 10'd084 }; 
        'd0540: dout <= { 2'd1, 8'd115, 10'd347 }; 
        'd0541: dout <= { 2'd1, 8'd044, 10'd332 }; 
        'd0542: dout <= { 2'd2, 8'd093, 10'd189 }; 
        'd0543: dout <= { 2'd1, 8'd095, 10'd121 }; 
        'd0544: dout <= { 2'd1, 8'd113, 10'd129 }; 
        'd0545: dout <= { 2'd2, 8'd082, 10'd013 }; 
        'd0546: dout <= { 2'd1, 8'd071, 10'd242 }; 
        'd0547: dout <= { 2'd1, 8'd101, 10'd308 }; 
        'd0548: dout <= { 2'd2, 8'd020, 10'd332 }; 
        'd0549: dout <= { 2'd1, 8'd099, 10'd079 }; 
        'd0550: dout <= { 2'd1, 8'd072, 10'd279 }; 
        'd0551: dout <= { 2'd2, 8'd033, 10'd005 }; 
        'd0552: dout <= { 2'd1, 8'd111, 10'd107 }; 
        'd0553: dout <= { 2'd1, 8'd017, 10'd176 }; 
        'd0554: dout <= { 2'd2, 8'd008, 10'd330 }; 
        'd0555: dout <= { 2'd1, 8'd084, 10'd318 }; 
        'd0556: dout <= { 2'd1, 8'd001, 10'd228 }; 
        'd0557: dout <= { 2'd2, 8'd017, 10'd245 }; 
        'd0558: dout <= { 2'd1, 8'd059, 10'd024 }; 
        'd0559: dout <= { 2'd1, 8'd092, 10'd084 }; 
        'd0560: dout <= { 2'd2, 8'd119, 10'd303 }; 
        'd0561: dout <= { 2'd1, 8'd054, 10'd242 }; 
        'd0562: dout <= { 2'd1, 8'd077, 10'd044 }; 
        'd0563: dout <= { 2'd2, 8'd024, 10'd160 }; 
        'd0564: dout <= { 2'd1, 8'd082, 10'd079 }; 
        'd0565: dout <= { 2'd1, 8'd076, 10'd203 }; 
        'd0566: dout <= { 2'd2, 8'd077, 10'd238 }; 
        'd0567: dout <= { 2'd1, 8'd097, 10'd334 }; 
        'd0568: dout <= { 2'd1, 8'd046, 10'd019 }; 
        'd0569: dout <= { 2'd2, 8'd064, 10'd112 }; 
        'd0570: dout <= { 2'd1, 8'd114, 10'd056 }; 
        'd0571: dout <= { 2'd1, 8'd103, 10'd179 }; 
        'd0572: dout <= { 2'd2, 8'd036, 10'd354 }; 
        'd0573: dout <= { 2'd1, 8'd091, 10'd338 }; 
        'd0574: dout <= { 2'd1, 8'd090, 10'd356 }; 
        'd0575: dout <= { 2'd2, 8'd029, 10'd214 }; 
        'd0576: dout <= { 2'd1, 8'd117, 10'd262 }; 
        'd0577: dout <= { 2'd1, 8'd098, 10'd267 }; 
        'd0578: dout <= { 2'd2, 8'd102, 10'd317 }; 
        'd0579: dout <= { 2'd1, 8'd024, 10'd155 }; 
        'd0580: dout <= { 2'd1, 8'd107, 10'd348 }; 
        'd0581: dout <= { 2'd2, 8'd056, 10'd327 }; 
        'd0582: dout <= { 2'd1, 8'd000, 10'd313 }; 
        'd0583: dout <= { 2'd1, 8'd015, 10'd119 }; 
        'd0584: dout <= { 2'd2, 8'd045, 10'd135 }; 
        'd0585: dout <= { 2'd1, 8'd101, 10'd056 }; 
        'd0586: dout <= { 2'd1, 8'd079, 10'd180 }; 
        'd0587: dout <= { 2'd2, 8'd010, 10'd263 }; 
        'd0588: dout <= { 2'd1, 8'd019, 10'd211 }; 
        'd0589: dout <= { 2'd1, 8'd003, 10'd209 }; 
        'd0590: dout <= { 2'd2, 8'd001, 10'd184 }; 
        'd0591: dout <= { 2'd1, 8'd007, 10'd067 }; 
        'd0592: dout <= { 2'd1, 8'd097, 10'd005 }; 
        'd0593: dout <= { 2'd2, 8'd108, 10'd293 }; 
        'd0594: dout <= { 2'd1, 8'd044, 10'd082 }; 
        'd0595: dout <= { 2'd1, 8'd033, 10'd142 }; 
        'd0596: dout <= { 2'd2, 8'd075, 10'd166 }; 
        'd0597: dout <= { 2'd1, 8'd088, 10'd223 }; 
        'd0598: dout <= { 2'd1, 8'd085, 10'd293 }; 
        'd0599: dout <= { 2'd2, 8'd110, 10'd069 }; 
        'd0600: dout <= { 2'd1, 8'd058, 10'd155 }; 
        'd0601: dout <= { 2'd1, 8'd054, 10'd134 }; 
        'd0602: dout <= { 2'd2, 8'd047, 10'd123 }; 
        'd0603: dout <= { 2'd1, 8'd081, 10'd101 }; 
        'd0604: dout <= { 2'd1, 8'd064, 10'd274 }; 
        'd0605: dout <= { 2'd2, 8'd115, 10'd041 }; 
        'd0606: dout <= { 2'd1, 8'd036, 10'd210 }; 
        'd0607: dout <= { 2'd1, 8'd016, 10'd010 }; 
        'd0608: dout <= { 2'd2, 8'd106, 10'd324 }; 
        'd0609: dout <= { 2'd1, 8'd034, 10'd358 }; 
        'd0610: dout <= { 2'd1, 8'd062, 10'd206 }; 
        'd0611: dout <= { 2'd2, 8'd041, 10'd072 }; 
        'd0612: dout <= { 2'd1, 8'd001, 10'd236 }; 
        'd0613: dout <= { 2'd1, 8'd012, 10'd041 }; 
        'd0614: dout <= { 2'd2, 8'd049, 10'd285 }; 
        'd0615: dout <= { 2'd1, 8'd027, 10'd034 }; 
        'd0616: dout <= { 2'd1, 8'd102, 10'd244 }; 
        'd0617: dout <= { 2'd2, 8'd084, 10'd267 }; 
        'd0618: dout <= { 2'd1, 8'd077, 10'd184 }; 
        'd0619: dout <= { 2'd1, 8'd104, 10'd021 }; 
        'd0620: dout <= { 2'd2, 8'd068, 10'd120 }; 
        'd0621: dout <= { 2'd1, 8'd028, 10'd323 }; 
        'd0622: dout <= { 2'd1, 8'd081, 10'd225 }; 
        'd0623: dout <= { 2'd2, 8'd016, 10'd066 }; 
        'd0624: dout <= { 2'd1, 8'd048, 10'd036 }; 
        'd0625: dout <= { 2'd1, 8'd108, 10'd217 }; 
        'd0626: dout <= { 2'd2, 8'd018, 10'd088 }; 
        'd0627: dout <= { 2'd1, 8'd033, 10'd211 }; 
        'd0628: dout <= { 2'd1, 8'd042, 10'd034 }; 
        'd0629: dout <= { 2'd3, 8'd031, 10'd331 }; 
        // Q=108, BaseAddr=630
        'd0630: dout <= { 2'd1, 8'd093, 10'd290 }; 
        'd0631: dout <= { 2'd1, 8'd042, 10'd174 }; 
        'd0632: dout <= { 2'd1, 8'd048, 10'd267 }; 
        'd0633: dout <= { 2'd1, 8'd083, 10'd008 }; 
        'd0634: dout <= { 2'd1, 8'd046, 10'd213 }; 
        'd0635: dout <= { 2'd1, 8'd012, 10'd134 }; 
        'd0636: dout <= { 2'd1, 8'd013, 10'd137 }; 
        'd0637: dout <= { 2'd1, 8'd000, 10'd046 }; 
        'd0638: dout <= { 2'd1, 8'd023, 10'd004 }; 
        'd0639: dout <= { 2'd1, 8'd071, 10'd311 }; 
        'd0640: dout <= { 2'd1, 8'd034, 10'd154 }; 
        'd0641: dout <= { 2'd2, 8'd000, 10'd176 }; 
        'd0642: dout <= { 2'd1, 8'd104, 10'd121 }; 
        'd0643: dout <= { 2'd1, 8'd067, 10'd184 }; 
        'd0644: dout <= { 2'd1, 8'd070, 10'd123 }; 
        'd0645: dout <= { 2'd1, 8'd003, 10'd127 }; 
        'd0646: dout <= { 2'd1, 8'd084, 10'd056 }; 
        'd0647: dout <= { 2'd1, 8'd106, 10'd185 }; 
        'd0648: dout <= { 2'd1, 8'd020, 10'd315 }; 
        'd0649: dout <= { 2'd1, 8'd050, 10'd124 }; 
        'd0650: dout <= { 2'd1, 8'd094, 10'd258 }; 
        'd0651: dout <= { 2'd1, 8'd073, 10'd155 }; 
        'd0652: dout <= { 2'd1, 8'd027, 10'd274 }; 
        'd0653: dout <= { 2'd2, 8'd029, 10'd153 }; 
        'd0654: dout <= { 2'd1, 8'd095, 10'd013 }; 
        'd0655: dout <= { 2'd1, 8'd107, 10'd296 }; 
        'd0656: dout <= { 2'd1, 8'd058, 10'd138 }; 
        'd0657: dout <= { 2'd1, 8'd022, 10'd107 }; 
        'd0658: dout <= { 2'd1, 8'd080, 10'd103 }; 
        'd0659: dout <= { 2'd1, 8'd037, 10'd085 }; 
        'd0660: dout <= { 2'd1, 8'd009, 10'd097 }; 
        'd0661: dout <= { 2'd1, 8'd058, 10'd213 }; 
        'd0662: dout <= { 2'd1, 8'd048, 10'd286 }; 
        'd0663: dout <= { 2'd1, 8'd072, 10'd165 }; 
        'd0664: dout <= { 2'd1, 8'd012, 10'd224 }; 
        'd0665: dout <= { 2'd2, 8'd045, 10'd230 }; 
        'd0666: dout <= { 2'd1, 8'd090, 10'd300 }; 
        'd0667: dout <= { 2'd1, 8'd050, 10'd167 }; 
        'd0668: dout <= { 2'd1, 8'd079, 10'd166 }; 
        'd0669: dout <= { 2'd1, 8'd097, 10'd045 }; 
        'd0670: dout <= { 2'd1, 8'd049, 10'd067 }; 
        'd0671: dout <= { 2'd1, 8'd105, 10'd296 }; 
        'd0672: dout <= { 2'd1, 8'd030, 10'd176 }; 
        'd0673: dout <= { 2'd1, 8'd024, 10'd066 }; 
        'd0674: dout <= { 2'd1, 8'd066, 10'd115 }; 
        'd0675: dout <= { 2'd1, 8'd091, 10'd124 }; 
        'd0676: dout <= { 2'd1, 8'd076, 10'd229 }; 
        'd0677: dout <= { 2'd2, 8'd051, 10'd201 }; 
        'd0678: dout <= { 2'd1, 8'd029, 10'd299 }; 
        'd0679: dout <= { 2'd1, 8'd039, 10'd100 }; 
        'd0680: dout <= { 2'd1, 8'd068, 10'd144 }; 
        'd0681: dout <= { 2'd1, 8'd041, 10'd310 }; 
        'd0682: dout <= { 2'd1, 8'd026, 10'd213 }; 
        'd0683: dout <= { 2'd1, 8'd062, 10'd098 }; 
        'd0684: dout <= { 2'd1, 8'd100, 10'd242 }; 
        'd0685: dout <= { 2'd1, 8'd088, 10'd182 }; 
        'd0686: dout <= { 2'd1, 8'd005, 10'd201 }; 
        'd0687: dout <= { 2'd1, 8'd064, 10'd340 }; 
        'd0688: dout <= { 2'd1, 8'd024, 10'd074 }; 
        'd0689: dout <= { 2'd2, 8'd017, 10'd119 }; 
        'd0690: dout <= { 2'd1, 8'd065, 10'd329 }; 
        'd0691: dout <= { 2'd1, 8'd005, 10'd103 }; 
        'd0692: dout <= { 2'd1, 8'd020, 10'd166 }; 
        'd0693: dout <= { 2'd1, 8'd024, 10'd242 }; 
        'd0694: dout <= { 2'd1, 8'd041, 10'd136 }; 
        'd0695: dout <= { 2'd1, 8'd083, 10'd295 }; 
        'd0696: dout <= { 2'd1, 8'd004, 10'd189 }; 
        'd0697: dout <= { 2'd1, 8'd064, 10'd092 }; 
        'd0698: dout <= { 2'd1, 8'd106, 10'd072 }; 
        'd0699: dout <= { 2'd1, 8'd060, 10'd290 }; 
        'd0700: dout <= { 2'd1, 8'd102, 10'd257 }; 
        'd0701: dout <= { 2'd2, 8'd092, 10'd308 }; 
        'd0702: dout <= { 2'd1, 8'd085, 10'd130 }; 
        'd0703: dout <= { 2'd1, 8'd035, 10'd112 }; 
        'd0704: dout <= { 2'd1, 8'd019, 10'd335 }; 
        'd0705: dout <= { 2'd1, 8'd062, 10'd037 }; 
        'd0706: dout <= { 2'd1, 8'd028, 10'd333 }; 
        'd0707: dout <= { 2'd1, 8'd090, 10'd338 }; 
        'd0708: dout <= { 2'd1, 8'd002, 10'd312 }; 
        'd0709: dout <= { 2'd1, 8'd031, 10'd143 }; 
        'd0710: dout <= { 2'd1, 8'd054, 10'd014 }; 
        'd0711: dout <= { 2'd1, 8'd030, 10'd171 }; 
        'd0712: dout <= { 2'd1, 8'd089, 10'd117 }; 
        'd0713: dout <= { 2'd2, 8'd047, 10'd065 }; 
        'd0714: dout <= { 2'd1, 8'd018, 10'd161 }; 
        'd0715: dout <= { 2'd1, 8'd056, 10'd077 }; 
        'd0716: dout <= { 2'd1, 8'd013, 10'd328 }; 
        'd0717: dout <= { 2'd1, 8'd080, 10'd026 }; 
        'd0718: dout <= { 2'd1, 8'd104, 10'd010 }; 
        'd0719: dout <= { 2'd1, 8'd044, 10'd278 }; 
        'd0720: dout <= { 2'd1, 8'd098, 10'd238 }; 
        'd0721: dout <= { 2'd1, 8'd040, 10'd102 }; 
        'd0722: dout <= { 2'd1, 8'd107, 10'd050 }; 
        'd0723: dout <= { 2'd1, 8'd069, 10'd243 }; 
        'd0724: dout <= { 2'd1, 8'd021, 10'd298 }; 
        'd0725: dout <= { 2'd2, 8'd080, 10'd344 }; 
        'd0726: dout <= { 2'd1, 8'd026, 10'd141 }; 
        'd0727: dout <= { 2'd1, 8'd073, 10'd049 }; 
        'd0728: dout <= { 2'd1, 8'd028, 10'd160 }; 
        'd0729: dout <= { 2'd1, 8'd055, 10'd208 }; 
        'd0730: dout <= { 2'd1, 8'd017, 10'd324 }; 
        'd0731: dout <= { 2'd1, 8'd070, 10'd006 }; 
        'd0732: dout <= { 2'd1, 8'd056, 10'd048 }; 
        'd0733: dout <= { 2'd1, 8'd038, 10'd155 }; 
        'd0734: dout <= { 2'd1, 8'd019, 10'd214 }; 
        'd0735: dout <= { 2'd1, 8'd008, 10'd223 }; 
        'd0736: dout <= { 2'd1, 8'd067, 10'd190 }; 
        'd0737: dout <= { 2'd2, 8'd013, 10'd309 }; 
        'd0738: dout <= { 2'd1, 8'd023, 10'd254 }; 
        'd0739: dout <= { 2'd1, 8'd106, 10'd162 }; 
        'd0740: dout <= { 2'd1, 8'd054, 10'd042 }; 
        'd0741: dout <= { 2'd1, 8'd059, 10'd201 }; 
        'd0742: dout <= { 2'd1, 8'd018, 10'd206 }; 
        'd0743: dout <= { 2'd1, 8'd033, 10'd253 }; 
        'd0744: dout <= { 2'd1, 8'd052, 10'd281 }; 
        'd0745: dout <= { 2'd1, 8'd092, 10'd080 }; 
        'd0746: dout <= { 2'd1, 8'd088, 10'd051 }; 
        'd0747: dout <= { 2'd1, 8'd036, 10'd028 }; 
        'd0748: dout <= { 2'd1, 8'd007, 10'd312 }; 
        'd0749: dout <= { 2'd2, 8'd032, 10'd033 }; 
        'd0750: dout <= { 2'd1, 8'd078, 10'd063 }; 
        'd0751: dout <= { 2'd1, 8'd009, 10'd008 }; 
        'd0752: dout <= { 2'd1, 8'd089, 10'd101 }; 
        'd0753: dout <= { 2'd1, 8'd006, 10'd229 }; 
        'd0754: dout <= { 2'd1, 8'd034, 10'd192 }; 
        'd0755: dout <= { 2'd1, 8'd023, 10'd093 }; 
        'd0756: dout <= { 2'd1, 8'd095, 10'd123 }; 
        'd0757: dout <= { 2'd1, 8'd085, 10'd253 }; 
        'd0758: dout <= { 2'd1, 8'd083, 10'd235 }; 
        'd0759: dout <= { 2'd1, 8'd081, 10'd024 }; 
        'd0760: dout <= { 2'd1, 8'd086, 10'd064 }; 
        'd0761: dout <= { 2'd2, 8'd058, 10'd290 }; 
        'd0762: dout <= { 2'd1, 8'd061, 10'd140 }; 
        'd0763: dout <= { 2'd1, 8'd037, 10'd126 }; 
        'd0764: dout <= { 2'd1, 8'd049, 10'd319 }; 
        'd0765: dout <= { 2'd1, 8'd045, 10'd031 }; 
        'd0766: dout <= { 2'd1, 8'd060, 10'd035 }; 
        'd0767: dout <= { 2'd1, 8'd019, 10'd326 }; 
        'd0768: dout <= { 2'd1, 8'd010, 10'd144 }; 
        'd0769: dout <= { 2'd1, 8'd071, 10'd218 }; 
        'd0770: dout <= { 2'd1, 8'd002, 10'd355 }; 
        'd0771: dout <= { 2'd1, 8'd043, 10'd112 }; 
        'd0772: dout <= { 2'd1, 8'd031, 10'd180 }; 
        'd0773: dout <= { 2'd2, 8'd039, 10'd143 }; 
        'd0774: dout <= { 2'd1, 8'd066, 10'd123 }; 
        'd0775: dout <= { 2'd1, 8'd011, 10'd062 }; 
        'd0776: dout <= { 2'd1, 8'd057, 10'd219 }; 
        'd0777: dout <= { 2'd1, 8'd052, 10'd344 }; 
        'd0778: dout <= { 2'd1, 8'd074, 10'd238 }; 
        'd0779: dout <= { 2'd1, 8'd022, 10'd195 }; 
        'd0780: dout <= { 2'd1, 8'd059, 10'd069 }; 
        'd0781: dout <= { 2'd1, 8'd008, 10'd135 }; 
        'd0782: dout <= { 2'd1, 8'd074, 10'd092 }; 
        'd0783: dout <= { 2'd1, 8'd038, 10'd202 }; 
        'd0784: dout <= { 2'd1, 8'd079, 10'd262 }; 
        'd0785: dout <= { 2'd2, 8'd003, 10'd311 }; 
        'd0786: dout <= { 2'd1, 8'd094, 10'd115 }; 
        'd0787: dout <= { 2'd1, 8'd051, 10'd043 }; 
        'd0788: dout <= { 2'd1, 8'd038, 10'd344 }; 
        'd0789: dout <= { 2'd1, 8'd103, 10'd197 }; 
        'd0790: dout <= { 2'd1, 8'd039, 10'd173 }; 
        'd0791: dout <= { 2'd1, 8'd078, 10'd053 }; 
        'd0792: dout <= { 2'd1, 8'd054, 10'd066 }; 
        'd0793: dout <= { 2'd1, 8'd045, 10'd023 }; 
        'd0794: dout <= { 2'd1, 8'd020, 10'd277 }; 
        'd0795: dout <= { 2'd1, 8'd004, 10'd332 }; 
        'd0796: dout <= { 2'd1, 8'd042, 10'd262 }; 
        'd0797: dout <= { 2'd2, 8'd035, 10'd100 }; 
        'd0798: dout <= { 2'd1, 8'd047, 10'd317 }; 
        'd0799: dout <= { 2'd1, 8'd014, 10'd237 }; 
        'd0800: dout <= { 2'd1, 8'd086, 10'd305 }; 
        'd0801: dout <= { 2'd1, 8'd021, 10'd287 }; 
        'd0802: dout <= { 2'd1, 8'd091, 10'd196 }; 
        'd0803: dout <= { 2'd1, 8'd005, 10'd020 }; 
        'd0804: dout <= { 2'd1, 8'd099, 10'd201 }; 
        'd0805: dout <= { 2'd1, 8'd102, 10'd347 }; 
        'd0806: dout <= { 2'd1, 8'd095, 10'd010 }; 
        'd0807: dout <= { 2'd1, 8'd078, 10'd154 }; 
        'd0808: dout <= { 2'd1, 8'd015, 10'd203 }; 
        'd0809: dout <= { 2'd2, 8'd061, 10'd285 }; 
        'd0810: dout <= { 2'd1, 8'd076, 10'd252 }; 
        'd0811: dout <= { 2'd1, 8'd034, 10'd312 }; 
        'd0812: dout <= { 2'd1, 8'd032, 10'd063 }; 
        'd0813: dout <= { 2'd1, 8'd016, 10'd245 }; 
        'd0814: dout <= { 2'd1, 8'd107, 10'd254 }; 
        'd0815: dout <= { 2'd1, 8'd036, 10'd331 }; 
        'd0816: dout <= { 2'd1, 8'd101, 10'd168 }; 
        'd0817: dout <= { 2'd1, 8'd086, 10'd151 }; 
        'd0818: dout <= { 2'd1, 8'd011, 10'd166 }; 
        'd0819: dout <= { 2'd1, 8'd090, 10'd213 }; 
        'd0820: dout <= { 2'd1, 8'd100, 10'd177 }; 
        'd0821: dout <= { 2'd2, 8'd044, 10'd161 }; 
        'd0822: dout <= { 2'd1, 8'd099, 10'd107 }; 
        'd0823: dout <= { 2'd1, 8'd027, 10'd057 }; 
        'd0824: dout <= { 2'd1, 8'd044, 10'd358 }; 
        'd0825: dout <= { 2'd1, 8'd004, 10'd263 }; 
        'd0826: dout <= { 2'd1, 8'd057, 10'd325 }; 
        'd0827: dout <= { 2'd1, 8'd025, 10'd158 }; 
        'd0828: dout <= { 2'd1, 8'd066, 10'd129 }; 
        'd0829: dout <= { 2'd1, 8'd065, 10'd333 }; 
        'd0830: dout <= { 2'd1, 8'd040, 10'd139 }; 
        'd0831: dout <= { 2'd1, 8'd093, 10'd153 }; 
        'd0832: dout <= { 2'd1, 8'd022, 10'd052 }; 
        'd0833: dout <= { 2'd2, 8'd068, 10'd337 }; 
        'd0834: dout <= { 2'd1, 8'd033, 10'd145 }; 
        'd0835: dout <= { 2'd1, 8'd087, 10'd267 }; 
        'd0836: dout <= { 2'd1, 8'd001, 10'd243 }; 
        'd0837: dout <= { 2'd1, 8'd036, 10'd087 }; 
        'd0838: dout <= { 2'd1, 8'd011, 10'd108 }; 
        'd0839: dout <= { 2'd1, 8'd016, 10'd238 }; 
        'd0840: dout <= { 2'd1, 8'd053, 10'd244 }; 
        'd0841: dout <= { 2'd1, 8'd006, 10'd054 }; 
        'd0842: dout <= { 2'd1, 8'd099, 10'd294 }; 
        'd0843: dout <= { 2'd1, 8'd006, 10'd249 }; 
        'd0844: dout <= { 2'd1, 8'd098, 10'd074 }; 
        'd0845: dout <= { 2'd2, 8'd101, 10'd342 }; 
        'd0846: dout <= { 2'd1, 8'd010, 10'd226 }; 
        'd0847: dout <= { 2'd1, 8'd043, 10'd255 }; 
        'd0848: dout <= { 2'd1, 8'd075, 10'd073 }; 
        'd0849: dout <= { 2'd1, 8'd030, 10'd329 }; 
        'd0850: dout <= { 2'd1, 8'd079, 10'd349 }; 
        'd0851: dout <= { 2'd1, 8'd072, 10'd164 }; 
        'd0852: dout <= { 2'd1, 8'd042, 10'd105 }; 
        'd0853: dout <= { 2'd1, 8'd032, 10'd103 }; 
        'd0854: dout <= { 2'd1, 8'd055, 10'd350 }; 
        'd0855: dout <= { 2'd1, 8'd053, 10'd065 }; 
        'd0856: dout <= { 2'd1, 8'd085, 10'd200 }; 
        'd0857: dout <= { 2'd2, 8'd063, 10'd319 }; 
        'd0858: dout <= { 2'd1, 8'd069, 10'd101 }; 
        'd0859: dout <= { 2'd1, 8'd025, 10'd126 }; 
        'd0860: dout <= { 2'd1, 8'd081, 10'd286 }; 
        'd0861: dout <= { 2'd1, 8'd064, 10'd069 }; 
        'd0862: dout <= { 2'd1, 8'd063, 10'd110 }; 
        'd0863: dout <= { 2'd1, 8'd055, 10'd168 }; 
        'd0864: dout <= { 2'd1, 8'd047, 10'd048 }; 
        'd0865: dout <= { 2'd1, 8'd001, 10'd128 }; 
        'd0866: dout <= { 2'd1, 8'd041, 10'd181 }; 
        'd0867: dout <= { 2'd1, 8'd009, 10'd219 }; 
        'd0868: dout <= { 2'd1, 8'd026, 10'd103 }; 
        'd0869: dout <= { 2'd2, 8'd070, 10'd329 }; 
        'd0870: dout <= { 2'd1, 8'd008, 10'd177 }; 
        'd0871: dout <= { 2'd1, 8'd102, 10'd284 }; 
        'd0872: dout <= { 2'd1, 8'd082, 10'd061 }; 
        'd0873: dout <= { 2'd1, 8'd084, 10'd345 }; 
        'd0874: dout <= { 2'd1, 8'd094, 10'd152 }; 
        'd0875: dout <= { 2'd1, 8'd073, 10'd243 }; 
        'd0876: dout <= { 2'd1, 8'd082, 10'd217 }; 
        'd0877: dout <= { 2'd1, 8'd061, 10'd212 }; 
        'd0878: dout <= { 2'd1, 8'd084, 10'd058 }; 
        'd0879: dout <= { 2'd1, 8'd049, 10'd315 }; 
        'd0880: dout <= { 2'd1, 8'd097, 10'd081 }; 
        'd0881: dout <= { 2'd2, 8'd087, 10'd186 }; 
        'd0882: dout <= { 2'd1, 8'd101, 10'd323 }; 
        'd0883: dout <= { 2'd1, 8'd077, 10'd133 }; 
        'd0884: dout <= { 2'd1, 8'd072, 10'd237 }; 
        'd0885: dout <= { 2'd1, 8'd012, 10'd038 }; 
        'd0886: dout <= { 2'd1, 8'd103, 10'd027 }; 
        'd0887: dout <= { 2'd1, 8'd097, 10'd194 }; 
        'd0888: dout <= { 2'd1, 8'd048, 10'd345 }; 
        'd0889: dout <= { 2'd1, 8'd035, 10'd227 }; 
        'd0890: dout <= { 2'd1, 8'd103, 10'd228 }; 
        'd0891: dout <= { 2'd1, 8'd016, 10'd186 }; 
        'd0892: dout <= { 2'd1, 8'd010, 10'd230 }; 
        'd0893: dout <= { 2'd2, 8'd018, 10'd112 }; 
        'd0894: dout <= { 2'd1, 8'd063, 10'd353 }; 
        'd0895: dout <= { 2'd1, 8'd015, 10'd264 }; 
        'd0896: dout <= { 2'd1, 8'd040, 10'd121 }; 
        'd0897: dout <= { 2'd1, 8'd053, 10'd129 }; 
        'd0898: dout <= { 2'd1, 8'd021, 10'd013 }; 
        'd0899: dout <= { 2'd1, 8'd093, 10'd198 }; 
        'd0900: dout <= { 2'd1, 8'd027, 10'd285 }; 
        'd0901: dout <= { 2'd1, 8'd081, 10'd079 }; 
        'd0902: dout <= { 2'd1, 8'd105, 10'd242 }; 
        'd0903: dout <= { 2'd1, 8'd104, 10'd308 }; 
        'd0904: dout <= { 2'd1, 8'd057, 10'd332 }; 
        'd0905: dout <= { 2'd2, 8'd077, 10'd300 }; 
        'd0906: dout <= { 2'd1, 8'd071, 10'd054 }; 
        'd0907: dout <= { 2'd1, 8'd046, 10'd318 }; 
        'd0908: dout <= { 2'd1, 8'd017, 10'd228 }; 
        'd0909: dout <= { 2'd1, 8'd096, 10'd245 }; 
        'd0910: dout <= { 2'd1, 8'd003, 10'd213 }; 
        'd0911: dout <= { 2'd1, 8'd089, 10'd252 }; 
        'd0912: dout <= { 2'd1, 8'd015, 10'd354 }; 
        'd0913: dout <= { 2'd1, 8'd029, 10'd024 }; 
        'd0914: dout <= { 2'd1, 8'd050, 10'd084 }; 
        'd0915: dout <= { 2'd1, 8'd082, 10'd303 }; 
        'd0916: dout <= { 2'd1, 8'd062, 10'd199 }; 
        'd0917: dout <= { 2'd2, 8'd001, 10'd173 }; 
        'd0918: dout <= { 2'd1, 8'd007, 10'd160 }; 
        'd0919: dout <= { 2'd1, 8'd076, 10'd252 }; 
        'd0920: dout <= { 2'd2, 8'd025, 10'd176 }; 
        'd0921: dout <= { 2'd1, 8'd092, 10'd238 }; 
        'd0922: dout <= { 2'd1, 8'd043, 10'd294 }; 
        'd0923: dout <= { 2'd2, 8'd056, 10'd112 }; 
        'd0924: dout <= { 2'd1, 8'd088, 10'd112 }; 
        'd0925: dout <= { 2'd1, 8'd096, 10'd324 }; 
        'd0926: dout <= { 2'd2, 8'd014, 10'd289 }; 
        'd0927: dout <= { 2'd1, 8'd031, 10'd354 }; 
        'd0928: dout <= { 2'd1, 8'd014, 10'd309 }; 
        'd0929: dout <= { 2'd2, 8'd052, 10'd230 }; 
        'd0930: dout <= { 2'd1, 8'd002, 10'd214 }; 
        'd0931: dout <= { 2'd1, 8'd087, 10'd351 }; 
        'd0932: dout <= { 2'd2, 8'd096, 10'd275 }; 
        'd0933: dout <= { 2'd1, 8'd100, 10'd317 }; 
        'd0934: dout <= { 2'd1, 8'd075, 10'd097 }; 
        'd0935: dout <= { 2'd2, 8'd065, 10'd335 }; 
        'd0936: dout <= { 2'd1, 8'd091, 10'd327 }; 
        'd0937: dout <= { 2'd1, 8'd067, 10'd001 }; 
        'd0938: dout <= { 2'd2, 8'd075, 10'd066 }; 
        'd0939: dout <= { 2'd1, 8'd074, 10'd135 }; 
        'd0940: dout <= { 2'd1, 8'd077, 10'd353 }; 
        'd0941: dout <= { 2'd2, 8'd033, 10'd209 }; 
        'd0942: dout <= { 2'd1, 8'd000, 10'd263 }; 
        'd0943: dout <= { 2'd1, 8'd007, 10'd061 }; 
        'd0944: dout <= { 2'd2, 8'd046, 10'd009 }; 
        'd0945: dout <= { 2'd1, 8'd060, 10'd184 }; 
        'd0946: dout <= { 2'd1, 8'd068, 10'd032 }; 
        'd0947: dout <= { 2'd2, 8'd037, 10'd271 }; 
        'd0948: dout <= { 2'd1, 8'd105, 10'd293 }; 
        'd0949: dout <= { 2'd1, 8'd051, 10'd187 }; 
        'd0950: dout <= { 2'd2, 8'd028, 10'd075 }; 
        'd0951: dout <= { 2'd1, 8'd098, 10'd166 }; 
        'd0952: dout <= { 2'd1, 8'd069, 10'd336 }; 
        'd0953: dout <= { 2'd2, 8'd059, 10'd247 }; 
        'd0954: dout <= { 2'd1, 8'd091, 10'd069 }; 
        'd0955: dout <= { 2'd1, 8'd067, 10'd275 }; 
        'd0956: dout <= { 2'd2, 8'd088, 10'd125 }; 
        'd0957: dout <= { 2'd1, 8'd049, 10'd123 }; 
        'd0958: dout <= { 2'd1, 8'd045, 10'd240 }; 
        'd0959: dout <= { 2'd2, 8'd039, 10'd078 }; 
        'd0960: dout <= { 2'd1, 8'd032, 10'd134 }; 
        'd0961: dout <= { 2'd1, 8'd076, 10'd340 }; 
        'd0962: dout <= { 2'd2, 8'd054, 10'd182 }; 
        'd0963: dout <= { 2'd1, 8'd100, 10'd041 }; 
        'd0964: dout <= { 2'd1, 8'd027, 10'd234 }; 
        'd0965: dout <= { 2'd2, 8'd082, 10'd067 }; 
        'd0966: dout <= { 2'd1, 8'd099, 10'd324 }; 
        'd0967: dout <= { 2'd1, 8'd062, 10'd236 }; 
        'd0968: dout <= { 2'd2, 8'd002, 10'd137 }; 
        'd0969: dout <= { 2'd1, 8'd048, 10'd072 }; 
        'd0970: dout <= { 2'd1, 8'd107, 10'd001 }; 
        'd0971: dout <= { 2'd2, 8'd060, 10'd011 }; 
        'd0972: dout <= { 2'd1, 8'd068, 10'd285 }; 
        'd0973: dout <= { 2'd1, 8'd070, 10'd049 }; 
        'd0974: dout <= { 2'd2, 8'd011, 10'd160 }; 
        'd0975: dout <= { 2'd1, 8'd096, 10'd267 }; 
        'd0976: dout <= { 2'd1, 8'd009, 10'd280 }; 
        'd0977: dout <= { 2'd2, 8'd073, 10'd250 }; 
        'd0978: dout <= { 2'd1, 8'd102, 10'd120 }; 
        'd0979: dout <= { 2'd1, 8'd051, 10'd019 }; 
        'd0980: dout <= { 2'd2, 8'd006, 10'd150 }; 
        'd0981: dout <= { 2'd1, 8'd001, 10'd066 }; 
        'd0982: dout <= { 2'd1, 8'd094, 10'd296 }; 
        'd0983: dout <= { 2'd2, 8'd064, 10'd181 }; 
        'd0984: dout <= { 2'd1, 8'd008, 10'd088 }; 
        'd0985: dout <= { 2'd1, 8'd012, 10'd203 }; 
        'd0986: dout <= { 2'd2, 8'd061, 10'd359 }; 
        'd0987: dout <= { 2'd1, 8'd101, 10'd331 }; 
        'd0988: dout <= { 2'd1, 8'd058, 10'd312 }; 
        'd0989: dout <= { 2'd2, 8'd014, 10'd217 }; 
        'd0990: dout <= { 2'd1, 8'd021, 10'd173 }; 
        'd0991: dout <= { 2'd1, 8'd036, 10'd265 }; 
        'd0992: dout <= { 2'd2, 8'd075, 10'd167 }; 
        'd0993: dout <= { 2'd1, 8'd069, 10'd210 }; 
        'd0994: dout <= { 2'd1, 8'd024, 10'd254 }; 
        'd0995: dout <= { 2'd2, 8'd003, 10'd298 }; 
        'd0996: dout <= { 2'd1, 8'd041, 10'd261 }; 
        'd0997: dout <= { 2'd1, 8'd040, 10'd293 }; 
        'd0998: dout <= { 2'd2, 8'd028, 10'd279 }; 
        'd0999: dout <= { 2'd1, 8'd065, 10'd141 }; 
        'd1000: dout <= { 2'd1, 8'd059, 10'd078 }; 
        'd1001: dout <= { 2'd2, 8'd030, 10'd259 }; 
        'd1002: dout <= { 2'd1, 8'd084, 10'd137 }; 
        'd1003: dout <= { 2'd1, 8'd050, 10'd123 }; 
        'd1004: dout <= { 2'd2, 8'd056, 10'd116 }; 
        'd1005: dout <= { 2'd1, 8'd026, 10'd265 }; 
        'd1006: dout <= { 2'd1, 8'd074, 10'd023 }; 
        'd1007: dout <= { 2'd2, 8'd031, 10'd182 }; 
        'd1008: dout <= { 2'd1, 8'd103, 10'd057 }; 
        'd1009: dout <= { 2'd1, 8'd071, 10'd041 }; 
        'd1010: dout <= { 2'd2, 8'd092, 10'd243 }; 
        'd1011: dout <= { 2'd1, 8'd072, 10'd110 }; 
        'd1012: dout <= { 2'd1, 8'd090, 10'd262 }; 
        'd1013: dout <= { 2'd2, 8'd089, 10'd077 }; 
        'd1014: dout <= { 2'd1, 8'd025, 10'd098 }; 
        'd1015: dout <= { 2'd1, 8'd097, 10'd008 }; 
        'd1016: dout <= { 2'd2, 8'd022, 10'd070 }; 
        'd1017: dout <= { 2'd1, 8'd055, 10'd096 }; 
        'd1018: dout <= { 2'd1, 8'd015, 10'd122 }; 
        'd1019: dout <= { 2'd2, 8'd034, 10'd248 }; 
        'd1020: dout <= { 2'd1, 8'd046, 10'd147 }; 
        'd1021: dout <= { 2'd1, 8'd042, 10'd339 }; 
        'd1022: dout <= { 2'd2, 8'd066, 10'd198 }; 
        'd1023: dout <= { 2'd1, 8'd016, 10'd097 }; 
        'd1024: dout <= { 2'd1, 8'd020, 10'd014 }; 
        'd1025: dout <= { 2'd2, 8'd017, 10'd011 }; 
        'd1026: dout <= { 2'd1, 8'd095, 10'd282 }; 
        'd1027: dout <= { 2'd1, 8'd086, 10'd337 }; 
        'd1028: dout <= { 2'd2, 8'd013, 10'd205 }; 
        'd1029: dout <= { 2'd1, 8'd080, 10'd047 }; 
        'd1030: dout <= { 2'd1, 8'd098, 10'd104 }; 
        'd1031: dout <= { 2'd2, 8'd007, 10'd317 }; 
        'd1032: dout <= { 2'd1, 8'd104, 10'd264 }; 
        'd1033: dout <= { 2'd1, 8'd053, 10'd327 }; 
        'd1034: dout <= { 2'd2, 8'd038, 10'd123 }; 
        'd1035: dout <= { 2'd1, 8'd106, 10'd082 }; 
        'd1036: dout <= { 2'd1, 8'd081, 10'd013 }; 
        'd1037: dout <= { 2'd2, 8'd018, 10'd196 }; 
        'd1038: dout <= { 2'd1, 8'd105, 10'd217 }; 
        'd1039: dout <= { 2'd1, 8'd057, 10'd161 }; 
        'd1040: dout <= { 2'd2, 8'd029, 10'd329 }; 
        'd1041: dout <= { 2'd1, 8'd085, 10'd306 }; 
        'd1042: dout <= { 2'd1, 8'd037, 10'd107 }; 
        'd1043: dout <= { 2'd2, 8'd023, 10'd184 }; 
        'd1044: dout <= { 2'd1, 8'd005, 10'd314 }; 
        'd1045: dout <= { 2'd1, 8'd087, 10'd072 }; 
        'd1046: dout <= { 2'd2, 8'd063, 10'd311 }; 
        'd1047: dout <= { 2'd1, 8'd083, 10'd185 }; 
        'd1048: dout <= { 2'd1, 8'd035, 10'd262 }; 
        'd1049: dout <= { 2'd2, 8'd010, 10'd099 }; 
        'd1050: dout <= { 2'd1, 8'd019, 10'd122 }; 
        'd1051: dout <= { 2'd1, 8'd047, 10'd195 }; 
        'd1052: dout <= { 2'd2, 8'd043, 10'd202 }; 
        'd1053: dout <= { 2'd1, 8'd044, 10'd040 }; 
        'd1054: dout <= { 2'd1, 8'd033, 10'd288 }; 
        'd1055: dout <= { 2'd2, 8'd052, 10'd044 }; 
        'd1056: dout <= { 2'd1, 8'd077, 10'd051 }; 
        'd1057: dout <= { 2'd1, 8'd093, 10'd018 }; 
        'd1058: dout <= { 2'd2, 8'd078, 10'd044 }; 
        'd1059: dout <= { 2'd1, 8'd000, 10'd284 }; 
        'd1060: dout <= { 2'd1, 8'd079, 10'd156 }; 
        'd1061: dout <= { 2'd3, 8'd004, 10'd137 }; 
        // Q=90, BaseAddr=1062
        'd1062: dout <= { 2'd1, 8'd054, 10'd000 }; 
        'd1063: dout <= { 2'd1, 8'd048, 10'd103 }; 
        'd1064: dout <= { 2'd1, 8'd082, 10'd159 }; 
        'd1065: dout <= { 2'd1, 8'd021, 10'd306 }; 
        'd1066: dout <= { 2'd1, 8'd089, 10'd298 }; 
        'd1067: dout <= { 2'd1, 8'd049, 10'd113 }; 
        'd1068: dout <= { 2'd1, 8'd014, 10'd028 }; 
        'd1069: dout <= { 2'd2, 8'd047, 10'd095 }; 
        'd1070: dout <= { 2'd1, 8'd055, 10'd000 }; 
        'd1071: dout <= { 2'd1, 8'd063, 10'd080 }; 
        'd1072: dout <= { 2'd1, 8'd045, 10'd051 }; 
        'd1073: dout <= { 2'd1, 8'd010, 10'd028 }; 
        'd1074: dout <= { 2'd1, 8'd050, 10'd312 }; 
        'd1075: dout <= { 2'd1, 8'd063, 10'd033 }; 
        'd1076: dout <= { 2'd1, 8'd070, 10'd264 }; 
        'd1077: dout <= { 2'd2, 8'd051, 10'd040 }; 
        'd1078: dout <= { 2'd1, 8'd056, 10'd000 }; 
        'd1079: dout <= { 2'd1, 8'd071, 10'd274 }; 
        'd1080: dout <= { 2'd1, 8'd003, 10'd262 }; 
        'd1081: dout <= { 2'd1, 8'd026, 10'd289 }; 
        'd1082: dout <= { 2'd1, 8'd019, 10'd192 }; 
        'd1083: dout <= { 2'd1, 8'd080, 10'd063 }; 
        'd1084: dout <= { 2'd1, 8'd072, 10'd008 }; 
        'd1085: dout <= { 2'd2, 8'd079, 10'd101 }; 
        'd1086: dout <= { 2'd1, 8'd057, 10'd000 }; 
        'd1087: dout <= { 2'd1, 8'd051, 10'd064 }; 
        'd1088: dout <= { 2'd1, 8'd054, 10'd290 }; 
        'd1089: dout <= { 2'd1, 8'd023, 10'd207 }; 
        'd1090: dout <= { 2'd1, 8'd031, 10'd128 }; 
        'd1091: dout <= { 2'd1, 8'd057, 10'd171 }; 
        'd1092: dout <= { 2'd1, 8'd005, 10'd152 }; 
        'd1093: dout <= { 2'd2, 8'd064, 10'd180 }; 
        'd1094: dout <= { 2'd1, 8'd058, 10'd000 }; 
        'd1095: dout <= { 2'd1, 8'd010, 10'd140 }; 
        'd1096: dout <= { 2'd1, 8'd007, 10'd126 }; 
        'd1097: dout <= { 2'd1, 8'd058, 10'd319 }; 
        'd1098: dout <= { 2'd1, 8'd002, 10'd031 }; 
        'd1099: dout <= { 2'd1, 8'd024, 10'd035 }; 
        'd1100: dout <= { 2'd1, 8'd031, 10'd326 }; 
        'd1101: dout <= { 2'd2, 8'd037, 10'd144 }; 
        'd1102: dout <= { 2'd1, 8'd059, 10'd000 }; 
        'd1103: dout <= { 2'd1, 8'd049, 10'd186 }; 
        'd1104: dout <= { 2'd1, 8'd088, 10'd177 }; 
        'd1105: dout <= { 2'd1, 8'd029, 10'd238 }; 
        'd1106: dout <= { 2'd1, 8'd045, 10'd068 }; 
        'd1107: dout <= { 2'd1, 8'd052, 10'd235 }; 
        'd1108: dout <= { 2'd1, 8'd010, 10'd176 }; 
        'd1109: dout <= { 2'd2, 8'd036, 10'd035 }; 
        'd1110: dout <= { 2'd1, 8'd060, 10'd000 }; 
        'd1111: dout <= { 2'd1, 8'd056, 10'd344 }; 
        'd1112: dout <= { 2'd1, 8'd029, 10'd238 }; 
        'd1113: dout <= { 2'd1, 8'd068, 10'd195 }; 
        'd1114: dout <= { 2'd1, 8'd003, 10'd069 }; 
        'd1115: dout <= { 2'd1, 8'd016, 10'd135 }; 
        'd1116: dout <= { 2'd1, 8'd054, 10'd092 }; 
        'd1117: dout <= { 2'd2, 8'd032, 10'd202 }; 
        'd1118: dout <= { 2'd1, 8'd061, 10'd000 }; 
        'd1119: dout <= { 2'd1, 8'd066, 10'd253 }; 
        'd1120: dout <= { 2'd1, 8'd083, 10'd157 }; 
        'd1121: dout <= { 2'd1, 8'd077, 10'd125 }; 
        'd1122: dout <= { 2'd1, 8'd046, 10'd065 }; 
        'd1123: dout <= { 2'd1, 8'd088, 10'd007 }; 
        'd1124: dout <= { 2'd1, 8'd027, 10'd130 }; 
        'd1125: dout <= { 2'd2, 8'd038, 10'd103 }; 
        'd1126: dout <= { 2'd1, 8'd062, 10'd000 }; 
        'd1127: dout <= { 2'd1, 8'd021, 10'd023 }; 
        'd1128: dout <= { 2'd1, 8'd011, 10'd277 }; 
        'd1129: dout <= { 2'd1, 8'd086, 10'd332 }; 
        'd1130: dout <= { 2'd1, 8'd054, 10'd262 }; 
        'd1131: dout <= { 2'd1, 8'd013, 10'd100 }; 
        'd1132: dout <= { 2'd1, 8'd017, 10'd173 }; 
        'd1133: dout <= { 2'd2, 8'd044, 10'd060 }; 
        'd1134: dout <= { 2'd1, 8'd063, 10'd000 }; 
        'd1135: dout <= { 2'd1, 8'd067, 10'd246 }; 
        'd1136: dout <= { 2'd1, 8'd023, 10'd044 }; 
        'd1137: dout <= { 2'd1, 8'd074, 10'd187 }; 
        'd1138: dout <= { 2'd1, 8'd004, 10'd317 }; 
        'd1139: dout <= { 2'd1, 8'd085, 10'd237 }; 
        'd1140: dout <= { 2'd1, 8'd074, 10'd305 }; 
        'd1141: dout <= { 2'd2, 8'd082, 10'd287 }; 
        'd1142: dout <= { 2'd1, 8'd064, 10'd000 }; 
        'd1143: dout <= { 2'd1, 8'd037, 10'd285 }; 
        'd1144: dout <= { 2'd1, 8'd001, 10'd050 }; 
        'd1145: dout <= { 2'd1, 8'd053, 10'd246 }; 
        'd1146: dout <= { 2'd1, 8'd085, 10'd162 }; 
        'd1147: dout <= { 2'd1, 8'd038, 10'd164 }; 
        'd1148: dout <= { 2'd1, 8'd048, 10'd179 }; 
        'd1149: dout <= { 2'd2, 8'd001, 10'd061 }; 
        'd1150: dout <= { 2'd1, 8'd065, 10'd000 }; 
        'd1151: dout <= { 2'd1, 8'd020, 10'd050 }; 
        'd1152: dout <= { 2'd1, 8'd084, 10'd189 }; 
        'd1153: dout <= { 2'd1, 8'd087, 10'd259 }; 
        'd1154: dout <= { 2'd1, 8'd034, 10'd047 }; 
        'd1155: dout <= { 2'd1, 8'd050, 10'd248 }; 
        'd1156: dout <= { 2'd1, 8'd021, 10'd188 }; 
        'd1157: dout <= { 2'd2, 8'd016, 10'd239 }; 
        'd1158: dout <= { 2'd1, 8'd066, 10'd000 }; 
        'd1159: dout <= { 2'd1, 8'd050, 10'd116 }; 
        'd1160: dout <= { 2'd1, 8'd062, 10'd068 }; 
        'd1161: dout <= { 2'd1, 8'd060, 10'd359 }; 
        'd1162: dout <= { 2'd1, 8'd057, 10'd106 }; 
        'd1163: dout <= { 2'd1, 8'd061, 10'd342 }; 
        'd1164: dout <= { 2'd1, 8'd034, 10'd288 }; 
        'd1165: dout <= { 2'd2, 8'd062, 10'd030 }; 
        'd1166: dout <= { 2'd1, 8'd067, 10'd000 }; 
        'd1167: dout <= { 2'd1, 8'd070, 10'd245 }; 
        'd1168: dout <= { 2'd1, 8'd005, 10'd254 }; 
        'd1169: dout <= { 2'd1, 8'd080, 10'd331 }; 
        'd1170: dout <= { 2'd1, 8'd027, 10'd168 }; 
        'd1171: dout <= { 2'd1, 8'd078, 10'd151 }; 
        'd1172: dout <= { 2'd1, 8'd015, 10'd166 }; 
        'd1173: dout <= { 2'd2, 8'd065, 10'd213 }; 
        'd1174: dout <= { 2'd1, 8'd068, 10'd000 }; 
        'd1175: dout <= { 2'd1, 8'd029, 10'd074 }; 
        'd1176: dout <= { 2'd1, 8'd048, 10'd204 }; 
        'd1177: dout <= { 2'd1, 8'd076, 10'd203 }; 
        'd1178: dout <= { 2'd1, 8'd018, 10'd110 }; 
        'd1179: dout <= { 2'd1, 8'd006, 10'd286 }; 
        'd1180: dout <= { 2'd1, 8'd043, 10'd060 }; 
        'd1181: dout <= { 2'd2, 8'd035, 10'd229 }; 
        'd1182: dout <= { 2'd1, 8'd069, 10'd000 }; 
        'd1183: dout <= { 2'd1, 8'd012, 10'd333 }; 
        'd1184: dout <= { 2'd1, 8'd019, 10'd139 }; 
        'd1185: dout <= { 2'd1, 8'd088, 10'd153 }; 
        'd1186: dout <= { 2'd1, 8'd066, 10'd052 }; 
        'd1187: dout <= { 2'd1, 8'd040, 10'd337 }; 
        'd1188: dout <= { 2'd1, 8'd033, 10'd111 }; 
        'd1189: dout <= { 2'd2, 8'd078, 10'd275 }; 
        'd1190: dout <= { 2'd1, 8'd070, 10'd000 }; 
        'd1191: dout <= { 2'd1, 8'd002, 10'd014 }; 
        'd1192: dout <= { 2'd1, 8'd042, 10'd311 }; 
        'd1193: dout <= { 2'd1, 8'd008, 10'd332 }; 
        'd1194: dout <= { 2'd1, 8'd013, 10'd145 }; 
        'd1195: dout <= { 2'd1, 8'd003, 10'd267 }; 
        'd1196: dout <= { 2'd1, 8'd081, 10'd243 }; 
        'd1197: dout <= { 2'd2, 8'd033, 10'd087 }; 
        'd1198: dout <= { 2'd1, 8'd071, 10'd000 }; 
        'd1199: dout <= { 2'd1, 8'd024, 10'd073 }; 
        'd1200: dout <= { 2'd1, 8'd032, 10'd329 }; 
        'd1201: dout <= { 2'd1, 8'd041, 10'd349 }; 
        'd1202: dout <= { 2'd1, 8'd071, 10'd164 }; 
        'd1203: dout <= { 2'd1, 8'd059, 10'd105 }; 
        'd1204: dout <= { 2'd1, 8'd065, 10'd103 }; 
        'd1205: dout <= { 2'd2, 8'd052, 10'd350 }; 
        'd1206: dout <= { 2'd1, 8'd072, 10'd000 }; 
        'd1207: dout <= { 2'd1, 8'd008, 10'd015 }; 
        'd1208: dout <= { 2'd1, 8'd064, 10'd071 }; 
        'd1209: dout <= { 2'd1, 8'd073, 10'd184 }; 
        'd1210: dout <= { 2'd1, 8'd014, 10'd226 }; 
        'd1211: dout <= { 2'd1, 8'd028, 10'd273 }; 
        'd1212: dout <= { 2'd1, 8'd084, 10'd006 }; 
        'd1213: dout <= { 2'd2, 8'd045, 10'd058 }; 
        'd1214: dout <= { 2'd1, 8'd073, 10'd000 }; 
        'd1215: dout <= { 2'd1, 8'd089, 10'd216 }; 
        'd1216: dout <= { 2'd1, 8'd025, 10'd003 }; 
        'd1217: dout <= { 2'd1, 8'd011, 10'd200 }; 
        'd1218: dout <= { 2'd1, 8'd020, 10'd034 }; 
        'd1219: dout <= { 2'd1, 8'd044, 10'd148 }; 
        'd1220: dout <= { 2'd1, 8'd022, 10'd089 }; 
        'd1221: dout <= { 2'd2, 8'd023, 10'd170 }; 
        'd1222: dout <= { 2'd1, 8'd074, 10'd000 }; 
        'd1223: dout <= { 2'd1, 8'd011, 10'd133 }; 
        'd1224: dout <= { 2'd1, 8'd070, 10'd016 }; 
        'd1225: dout <= { 2'd1, 8'd040, 10'd088 }; 
        'd1226: dout <= { 2'd1, 8'd042, 10'd238 }; 
        'd1227: dout <= { 2'd1, 8'd039, 10'd101 }; 
        'd1228: dout <= { 2'd1, 8'd030, 10'd126 }; 
        'd1229: dout <= { 2'd2, 8'd001, 10'd286 }; 
        'd1230: dout <= { 2'd1, 8'd075, 10'd000 }; 
        'd1231: dout <= { 2'd1, 8'd006, 10'd103 }; 
        'd1232: dout <= { 2'd1, 8'd046, 10'd329 }; 
        'd1233: dout <= { 2'd1, 8'd043, 10'd050 }; 
        'd1234: dout <= { 2'd1, 8'd009, 10'd341 }; 
        'd1235: dout <= { 2'd1, 8'd036, 10'd229 }; 
        'd1236: dout <= { 2'd1, 8'd051, 10'd243 }; 
        'd1237: dout <= { 2'd2, 8'd060, 10'd311 }; 
        'd1238: dout <= { 2'd1, 8'd076, 10'd000 }; 
        'd1239: dout <= { 2'd1, 8'd045, 10'd177 }; 
        'd1240: dout <= { 2'd1, 8'd074, 10'd284 }; 
        'd1241: dout <= { 2'd1, 8'd030, 10'd061 }; 
        'd1242: dout <= { 2'd1, 8'd069, 10'd345 }; 
        'd1243: dout <= { 2'd1, 8'd035, 10'd152 }; 
        'd1244: dout <= { 2'd1, 8'd079, 10'd243 }; 
        'd1245: dout <= { 2'd2, 8'd075, 10'd217 }; 
        'd1246: dout <= { 2'd1, 8'd077, 10'd000 }; 
        'd1247: dout <= { 2'd1, 8'd058, 10'd207 }; 
        'd1248: dout <= { 2'd1, 8'd018, 10'd051 }; 
        'd1249: dout <= { 2'd1, 8'd075, 10'd352 }; 
        'd1250: dout <= { 2'd1, 8'd015, 10'd335 }; 
        'd1251: dout <= { 2'd1, 8'd053, 10'd145 }; 
        'd1252: dout <= { 2'd1, 8'd086, 10'd118 }; 
        'd1253: dout <= { 2'd2, 8'd064, 10'd324 }; 
        'd1254: dout <= { 2'd1, 8'd078, 10'd000 }; 
        'd1255: dout <= { 2'd1, 8'd004, 10'd239 }; 
        'd1256: dout <= { 2'd1, 8'd077, 10'd256 }; 
        'd1257: dout <= { 2'd1, 8'd005, 10'd136 }; 
        'd1258: dout <= { 2'd1, 8'd025, 10'd289 }; 
        'd1259: dout <= { 2'd1, 8'd066, 10'd351 }; 
        'd1260: dout <= { 2'd1, 8'd071, 10'd284 }; 
        'd1261: dout <= { 2'd2, 8'd009, 10'd341 }; 
        'd1262: dout <= { 2'd1, 8'd079, 10'd000 }; 
        'd1263: dout <= { 2'd1, 8'd044, 10'd107 }; 
        'd1264: dout <= { 2'd1, 8'd036, 10'd277 }; 
        'd1265: dout <= { 2'd1, 8'd055, 10'd347 }; 
        'd1266: dout <= { 2'd1, 8'd028, 10'd332 }; 
        'd1267: dout <= { 2'd1, 8'd032, 10'd189 }; 
        'd1268: dout <= { 2'd1, 8'd018, 10'd273 }; 
        'd1269: dout <= { 2'd2, 8'd087, 10'd353 }; 
        'd1270: dout <= { 2'd1, 8'd080, 10'd000 }; 
        'd1271: dout <= { 2'd1, 8'd076, 10'd242 }; 
        'd1272: dout <= { 2'd1, 8'd057, 10'd308 }; 
        'd1273: dout <= { 2'd1, 8'd039, 10'd332 }; 
        'd1274: dout <= { 2'd1, 8'd000, 10'd300 }; 
        'd1275: dout <= { 2'd1, 8'd047, 10'd165 }; 
        'd1276: dout <= { 2'd1, 8'd069, 10'd126 }; 
        'd1277: dout <= { 2'd2, 8'd012, 10'd079 }; 
        'd1278: dout <= { 2'd1, 8'd081, 10'd000 }; 
        'd1279: dout <= { 2'd1, 8'd073, 10'd330 }; 
        'd1280: dout <= { 2'd1, 8'd000, 10'd259 }; 
        'd1281: dout <= { 2'd1, 8'd083, 10'd002 }; 
        'd1282: dout <= { 2'd1, 8'd017, 10'd054 }; 
        'd1283: dout <= { 2'd1, 8'd002, 10'd318 }; 
        'd1284: dout <= { 2'd1, 8'd025, 10'd228 }; 
        'd1285: dout <= { 2'd2, 8'd042, 10'd245 }; 
        'd1286: dout <= { 2'd1, 8'd082, 10'd000 }; 
        'd1287: dout <= { 2'd1, 8'd035, 10'd173 }; 
        'd1288: dout <= { 2'd1, 8'd071, 10'd062 }; 
        'd1289: dout <= { 2'd1, 8'd084, 10'd242 }; 
        'd1290: dout <= { 2'd1, 8'd007, 10'd044 }; 
        'd1291: dout <= { 2'd1, 8'd019, 10'd160 }; 
        'd1292: dout <= { 2'd1, 8'd077, 10'd252 }; 
        'd1293: dout <= { 2'd2, 8'd056, 10'd176 }; 
        'd1294: dout <= { 2'd1, 8'd083, 10'd000 }; 
        'd1295: dout <= { 2'd1, 8'd085, 10'd334 }; 
        'd1296: dout <= { 2'd1, 8'd049, 10'd019 }; 
        'd1297: dout <= { 2'd1, 8'd059, 10'd112 }; 
        'd1298: dout <= { 2'd1, 8'd063, 10'd324 }; 
        'd1299: dout <= { 2'd1, 8'd076, 10'd289 }; 
        'd1300: dout <= { 2'd1, 8'd026, 10'd117 }; 
        'd1301: dout <= { 2'd2, 8'd058, 10'd056 }; 
        'd1302: dout <= { 2'd1, 8'd084, 10'd000 }; 
        'd1303: dout <= { 2'd1, 8'd005, 10'd209 }; 
        'd1304: dout <= { 2'd1, 8'd015, 10'd184 }; 
        'd1305: dout <= { 2'd1, 8'd056, 10'd032 }; 
        'd1306: dout <= { 2'd1, 8'd067, 10'd271 }; 
        'd1307: dout <= { 2'd1, 8'd008, 10'd297 }; 
        'd1308: dout <= { 2'd1, 8'd000, 10'd067 }; 
        'd1309: dout <= { 2'd2, 8'd055, 10'd005 }; 
        'd1310: dout <= { 2'd1, 8'd085, 10'd000 }; 
        'd1311: dout <= { 2'd1, 8'd086, 10'd336 }; 
        'd1312: dout <= { 2'd1, 8'd068, 10'd247 }; 
        'd1313: dout <= { 2'd1, 8'd022, 10'd306 }; 
        'd1314: dout <= { 2'd1, 8'd061, 10'd223 }; 
        'd1315: dout <= { 2'd1, 8'd020, 10'd293 }; 
        'd1316: dout <= { 2'd1, 8'd037, 10'd069 }; 
        'd1317: dout <= { 2'd2, 8'd041, 10'd275 }; 
        'd1318: dout <= { 2'd1, 8'd086, 10'd000 }; 
        'd1319: dout <= { 2'd1, 8'd028, 10'd010 }; 
        'd1320: dout <= { 2'd1, 8'd086, 10'd324 }; 
        'd1321: dout <= { 2'd1, 8'd006, 10'd236 }; 
        'd1322: dout <= { 2'd1, 8'd070, 10'd137 }; 
        'd1323: dout <= { 2'd1, 8'd011, 10'd170 }; 
        'd1324: dout <= { 2'd1, 8'd089, 10'd358 }; 
        'd1325: dout <= { 2'd2, 8'd068, 10'd206 }; 
        'd1326: dout <= { 2'd1, 8'd087, 10'd000 }; 
        'd1327: dout <= { 2'd1, 8'd064, 10'd225 }; 
        'd1328: dout <= { 2'd1, 8'd085, 10'd066 }; 
        'd1329: dout <= { 2'd1, 8'd049, 10'd296 }; 
        'd1330: dout <= { 2'd1, 8'd012, 10'd181 }; 
        'd1331: dout <= { 2'd1, 8'd046, 10'd025 }; 
        'd1332: dout <= { 2'd1, 8'd004, 10'd036 }; 
        'd1333: dout <= { 2'd2, 8'd083, 10'd217 }; 
        'd1334: dout <= { 2'd1, 8'd088, 10'd000 }; 
        'd1335: dout <= { 2'd1, 8'd027, 10'd069 }; 
        'd1336: dout <= { 2'd1, 8'd063, 10'd132 }; 
        'd1337: dout <= { 2'd1, 8'd081, 10'd253 }; 
        'd1338: dout <= { 2'd1, 8'd072, 10'd173 }; 
        'd1339: dout <= { 2'd1, 8'd007, 10'd265 }; 
        'd1340: dout <= { 2'd1, 8'd082, 10'd167 }; 
        'd1341: dout <= { 2'd2, 8'd067, 10'd232 }; 
        'd1342: dout <= { 2'd1, 8'd089, 10'd000 }; 
        'd1343: dout <= { 2'd1, 8'd033, 10'd293 }; 
        'd1344: dout <= { 2'd1, 8'd058, 10'd279 }; 
        'd1345: dout <= { 2'd1, 8'd048, 10'd211 }; 
        'd1346: dout <= { 2'd1, 8'd024, 10'd204 }; 
        'd1347: dout <= { 2'd1, 8'd062, 10'd098 }; 
        'd1348: dout <= { 2'd1, 8'd029, 10'd141 }; 
        'd1349: dout <= { 2'd2, 8'd073, 10'd078 }; 
        'd1350: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd1351: dout <= { 2'd1, 8'd077, 10'd161 }; 
        'd1352: dout <= { 2'd2, 8'd035, 10'd277 }; 
        'd1353: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd1354: dout <= { 2'd1, 8'd038, 10'd043 }; 
        'd1355: dout <= { 2'd2, 8'd010, 10'd001 }; 
        'd1356: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd1357: dout <= { 2'd1, 8'd019, 10'd114 }; 
        'd1358: dout <= { 2'd2, 8'd060, 10'd002 }; 
        'd1359: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd1360: dout <= { 2'd1, 8'd072, 10'd267 }; 
        'd1361: dout <= { 2'd2, 8'd044, 10'd008 }; 
        'd1362: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd1363: dout <= { 2'd1, 8'd053, 10'd137 }; 
        'd1364: dout <= { 2'd2, 8'd033, 10'd046 }; 
        'd1365: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd1366: dout <= { 2'd1, 8'd001, 10'd154 }; 
        'd1367: dout <= { 2'd2, 8'd078, 10'd176 }; 
        'd1368: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd1369: dout <= { 2'd1, 8'd087, 10'd236 }; 
        'd1370: dout <= { 2'd2, 8'd056, 10'd011 }; 
        'd1371: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd1372: dout <= { 2'd1, 8'd068, 10'd058 }; 
        'd1373: dout <= { 2'd2, 8'd089, 10'd161 }; 
        'd1374: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd1375: dout <= { 2'd1, 8'd078, 10'd312 }; 
        'd1376: dout <= { 2'd2, 8'd059, 10'd089 }; 
        'd1377: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd1378: dout <= { 2'd1, 8'd023, 10'd184 }; 
        'd1379: dout <= { 2'd2, 8'd028, 10'd123 }; 
        'd1380: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd1381: dout <= { 2'd1, 8'd031, 10'd185 }; 
        'd1382: dout <= { 2'd2, 8'd013, 10'd315 }; 
        'd1383: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd1384: dout <= { 2'd1, 8'd030, 10'd155 }; 
        'd1385: dout <= { 2'd2, 8'd065, 10'd274 }; 
        'd1386: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd1387: dout <= { 2'd1, 8'd039, 10'd357 }; 
        'd1388: dout <= { 2'd2, 8'd079, 10'd199 }; 
        'd1389: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd1390: dout <= { 2'd1, 8'd017, 10'd121 }; 
        'd1391: dout <= { 2'd2, 8'd067, 10'd030 }; 
        'd1392: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd1393: dout <= { 2'd1, 8'd047, 10'd239 }; 
        'd1394: dout <= { 2'd2, 8'd038, 10'd042 }; 
        'd1395: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd1396: dout <= { 2'd1, 8'd036, 10'd296 }; 
        'd1397: dout <= { 2'd2, 8'd002, 10'd138 }; 
        'd1398: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd1399: dout <= { 2'd1, 8'd026, 10'd085 }; 
        'd1400: dout <= { 2'd2, 8'd024, 10'd097 }; 
        'd1401: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd1402: dout <= { 2'd1, 8'd055, 10'd165 }; 
        'd1403: dout <= { 2'd2, 8'd072, 10'd224 }; 
        'd1404: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd1405: dout <= { 2'd1, 8'd059, 10'd174 }; 
        'd1406: dout <= { 2'd2, 8'd076, 10'd273 }; 
        'd1407: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd1408: dout <= { 2'd1, 8'd082, 10'd354 }; 
        'd1409: dout <= { 2'd2, 8'd039, 10'd095 }; 
        'd1410: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd1411: dout <= { 2'd1, 8'd088, 10'd221 }; 
        'd1412: dout <= { 2'd2, 8'd017, 10'd302 }; 
        'd1413: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd1414: dout <= { 2'd1, 8'd060, 10'd300 }; 
        'd1415: dout <= { 2'd2, 8'd041, 10'd167 }; 
        'd1416: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd1417: dout <= { 2'd1, 8'd041, 10'd067 }; 
        'd1418: dout <= { 2'd2, 8'd009, 10'd296 }; 
        'd1419: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd1420: dout <= { 2'd1, 8'd043, 10'd115 }; 
        'd1421: dout <= { 2'd2, 8'd016, 10'd124 }; 
        'd1422: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd1423: dout <= { 2'd1, 8'd057, 10'd106 }; 
        'd1424: dout <= { 2'd2, 8'd050, 10'd148 }; 
        'd1425: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd1426: dout <= { 2'd1, 8'd061, 10'd078 }; 
        'd1427: dout <= { 2'd2, 8'd037, 10'd196 }; 
        'd1428: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd1429: dout <= { 2'd1, 8'd083, 10'd015 }; 
        'd1430: dout <= { 2'd2, 8'd073, 10'd216 }; 
        'd1431: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd1432: dout <= { 2'd1, 8'd015, 10'd299 }; 
        'd1433: dout <= { 2'd2, 8'd014, 10'd100 }; 
        'd1434: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd1435: dout <= { 2'd1, 8'd032, 10'd213 }; 
        'd1436: dout <= { 2'd2, 8'd080, 10'd098 }; 
        'd1437: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd1438: dout <= { 2'd1, 8'd062, 10'd201 }; 
        'd1439: dout <= { 2'd2, 8'd047, 10'd340 }; 
        'd1440: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd1441: dout <= { 2'd1, 8'd013, 10'd231 }; 
        'd1442: dout <= { 2'd2, 8'd027, 10'd019 }; 
        'd1443: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd1444: dout <= { 2'd1, 8'd014, 10'd131 }; 
        'd1445: dout <= { 2'd2, 8'd021, 10'd280 }; 
        'd1446: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd1447: dout <= { 2'd1, 8'd003, 10'd352 }; 
        'd1448: dout <= { 2'd2, 8'd053, 10'd197 }; 
        'd1449: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd1450: dout <= { 2'd1, 8'd084, 10'd329 }; 
        'd1451: dout <= { 2'd2, 8'd075, 10'd103 }; 
        'd1452: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd1453: dout <= { 2'd1, 8'd040, 10'd136 }; 
        'd1454: dout <= { 2'd2, 8'd061, 10'd295 }; 
        'd1455: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd1456: dout <= { 2'd1, 8'd046, 10'd072 }; 
        'd1457: dout <= { 2'd2, 8'd022, 10'd290 }; 
        'd1458: dout <= { 2'd1, 8'd036, 10'd000 }; 
        'd1459: dout <= { 2'd1, 8'd065, 10'd290 }; 
        'd1460: dout <= { 2'd2, 8'd081, 10'd124 }; 
        'd1461: dout <= { 2'd1, 8'd037, 10'd000 }; 
        'd1462: dout <= { 2'd1, 8'd016, 10'd085 }; 
        'd1463: dout <= { 2'd2, 8'd052, 10'd299 }; 
        'd1464: dout <= { 2'd1, 8'd038, 10'd000 }; 
        'd1465: dout <= { 2'd1, 8'd000, 10'd181 }; 
        'd1466: dout <= { 2'd2, 8'd020, 10'd094 }; 
        'd1467: dout <= { 2'd1, 8'd039, 10'd000 }; 
        'd1468: dout <= { 2'd1, 8'd074, 10'd130 }; 
        'd1469: dout <= { 2'd2, 8'd040, 10'd112 }; 
        'd1470: dout <= { 2'd1, 8'd040, 10'd000 }; 
        'd1471: dout <= { 2'd1, 8'd081, 10'd333 }; 
        'd1472: dout <= { 2'd2, 8'd006, 10'd338 }; 
        'd1473: dout <= { 2'd1, 8'd041, 10'd000 }; 
        'd1474: dout <= { 2'd1, 8'd075, 10'd014 }; 
        'd1475: dout <= { 2'd2, 8'd034, 10'd171 }; 
        'd1476: dout <= { 2'd1, 8'd042, 10'd000 }; 
        'd1477: dout <= { 2'd1, 8'd025, 10'd076 }; 
        'd1478: dout <= { 2'd2, 8'd012, 10'd197 }; 
        'd1479: dout <= { 2'd1, 8'd043, 10'd000 }; 
        'd1480: dout <= { 2'd1, 8'd009, 10'd353 }; 
        'd1481: dout <= { 2'd2, 8'd069, 10'd138 }; 
        'd1482: dout <= { 2'd1, 8'd044, 10'd000 }; 
        'd1483: dout <= { 2'd1, 8'd080, 10'd356 }; 
        'd1484: dout <= { 2'd2, 8'd031, 10'd233 }; 
        'd1485: dout <= { 2'd1, 8'd045, 10'd000 }; 
        'd1486: dout <= { 2'd1, 8'd018, 10'd161 }; 
        'd1487: dout <= { 2'd2, 8'd066, 10'd077 }; 
        'd1488: dout <= { 2'd1, 8'd046, 10'd000 }; 
        'd1489: dout <= { 2'd1, 8'd079, 10'd010 }; 
        'd1490: dout <= { 2'd2, 8'd004, 10'd278 }; 
        'd1491: dout <= { 2'd1, 8'd047, 10'd000 }; 
        'd1492: dout <= { 2'd1, 8'd054, 10'd050 }; 
        'd1493: dout <= { 2'd2, 8'd026, 10'd243 }; 
        'd1494: dout <= { 2'd1, 8'd048, 10'd000 }; 
        'd1495: dout <= { 2'd1, 8'd069, 10'd088 }; 
        'd1496: dout <= { 2'd2, 8'd087, 10'd241 }; 
        'd1497: dout <= { 2'd1, 8'd049, 10'd000 }; 
        'd1498: dout <= { 2'd1, 8'd022, 10'd055 }; 
        'd1499: dout <= { 2'd2, 8'd051, 10'd229 }; 
        'd1500: dout <= { 2'd1, 8'd050, 10'd000 }; 
        'd1501: dout <= { 2'd1, 8'd042, 10'd073 }; 
        'd1502: dout <= { 2'd2, 8'd030, 10'd030 }; 
        'd1503: dout <= { 2'd1, 8'd051, 10'd000 }; 
        'd1504: dout <= { 2'd1, 8'd052, 10'd141 }; 
        'd1505: dout <= { 2'd2, 8'd008, 10'd049 }; 
        'd1506: dout <= { 2'd1, 8'd052, 10'd000 }; 
        'd1507: dout <= { 2'd1, 8'd034, 10'd324 }; 
        'd1508: dout <= { 2'd2, 8'd055, 10'd006 }; 
        'd1509: dout <= { 2'd1, 8'd053, 10'd000 }; 
        'd1510: dout <= { 2'd1, 8'd007, 10'd214 }; 
        'd1511: dout <= { 2'd3, 8'd043, 10'd223 }; 
        // Q=72, BaseAddr=1512
        'd1512: dout <= { 2'd1, 8'd030, 10'd311 }; 
        'd1513: dout <= { 2'd1, 8'd058, 10'd142 }; 
        'd1514: dout <= { 2'd1, 8'd034, 10'd161 }; 
        'd1515: dout <= { 2'd1, 8'd053, 10'd277 }; 
        'd1516: dout <= { 2'd1, 8'd001, 10'd155 }; 
        'd1517: dout <= { 2'd1, 8'd042, 10'd040 }; 
        'd1518: dout <= { 2'd1, 8'd026, 10'd043 }; 
        'd1519: dout <= { 2'd1, 8'd027, 10'd001 }; 
        'd1520: dout <= { 2'd1, 8'd009, 10'd078 }; 
        'd1521: dout <= { 2'd1, 8'd000, 10'd237 }; 
        'd1522: dout <= { 2'd1, 8'd062, 10'd114 }; 
        'd1523: dout <= { 2'd2, 8'd035, 10'd002 }; 
        'd1524: dout <= { 2'd1, 8'd031, 10'd348 }; 
        'd1525: dout <= { 2'd1, 8'd018, 10'd225 }; 
        'd1526: dout <= { 2'd1, 8'd023, 10'd236 }; 
        'd1527: dout <= { 2'd1, 8'd036, 10'd011 }; 
        'd1528: dout <= { 2'd1, 8'd025, 10'd278 }; 
        'd1529: dout <= { 2'd1, 8'd024, 10'd356 }; 
        'd1530: dout <= { 2'd1, 8'd010, 10'd058 }; 
        'd1531: dout <= { 2'd1, 8'd037, 10'd161 }; 
        'd1532: dout <= { 2'd1, 8'd063, 10'd313 }; 
        'd1533: dout <= { 2'd1, 8'd025, 10'd240 }; 
        'd1534: dout <= { 2'd1, 8'd051, 10'd312 }; 
        'd1535: dout <= { 2'd2, 8'd055, 10'd089 }; 
        'd1536: dout <= { 2'd1, 8'd033, 10'd153 }; 
        'd1537: dout <= { 2'd1, 8'd029, 10'd317 }; 
        'd1538: dout <= { 2'd1, 8'd002, 10'd357 }; 
        'd1539: dout <= { 2'd1, 8'd060, 10'd199 }; 
        'd1540: dout <= { 2'd1, 8'd028, 10'd076 }; 
        'd1541: dout <= { 2'd1, 8'd021, 10'd267 }; 
        'd1542: dout <= { 2'd1, 8'd020, 10'd121 }; 
        'd1543: dout <= { 2'd1, 8'd017, 10'd030 }; 
        'd1544: dout <= { 2'd1, 8'd019, 10'd188 }; 
        'd1545: dout <= { 2'd1, 8'd042, 10'd157 }; 
        'd1546: dout <= { 2'd1, 8'd057, 10'd239 }; 
        'd1547: dout <= { 2'd2, 8'd045, 10'd042 }; 
        'd1548: dout <= { 2'd1, 8'd021, 10'd230 }; 
        'd1549: dout <= { 2'd1, 8'd049, 10'd308 }; 
        'd1550: dout <= { 2'd1, 8'd035, 10'd174 }; 
        'd1551: dout <= { 2'd1, 8'd061, 10'd273 }; 
        'd1552: dout <= { 2'd1, 8'd033, 10'd327 }; 
        'd1553: dout <= { 2'd1, 8'd035, 10'd160 }; 
        'd1554: dout <= { 2'd1, 8'd008, 10'd354 }; 
        'd1555: dout <= { 2'd1, 8'd013, 10'd095 }; 
        'd1556: dout <= { 2'd1, 8'd059, 10'd352 }; 
        'd1557: dout <= { 2'd1, 8'd034, 10'd072 }; 
        'd1558: dout <= { 2'd1, 8'd013, 10'd221 }; 
        'd1559: dout <= { 2'd2, 8'd022, 10'd302 }; 
        'd1560: dout <= { 2'd1, 8'd041, 10'd229 }; 
        'd1561: dout <= { 2'd1, 8'd015, 10'd201 }; 
        'd1562: dout <= { 2'd1, 8'd011, 10'd106 }; 
        'd1563: dout <= { 2'd1, 8'd059, 10'd148 }; 
        'd1564: dout <= { 2'd1, 8'd018, 10'd242 }; 
        'd1565: dout <= { 2'd1, 8'd031, 10'd154 }; 
        'd1566: dout <= { 2'd1, 8'd063, 10'd078 }; 
        'd1567: dout <= { 2'd1, 8'd043, 10'd196 }; 
        'd1568: dout <= { 2'd1, 8'd021, 10'd336 }; 
        'd1569: dout <= { 2'd1, 8'd048, 10'd291 }; 
        'd1570: dout <= { 2'd1, 8'd036, 10'd015 }; 
        'd1571: dout <= { 2'd2, 8'd068, 10'd216 }; 
        'd1572: dout <= { 2'd1, 8'd012, 10'd074 }; 
        'd1573: dout <= { 2'd1, 8'd068, 10'd119 }; 
        'd1574: dout <= { 2'd1, 8'd061, 10'd231 }; 
        'd1575: dout <= { 2'd1, 8'd066, 10'd019 }; 
        'd1576: dout <= { 2'd1, 8'd019, 10'd078 }; 
        'd1577: dout <= { 2'd1, 8'd036, 10'd090 }; 
        'd1578: dout <= { 2'd1, 8'd050, 10'd131 }; 
        'd1579: dout <= { 2'd1, 8'd029, 10'd280 }; 
        'd1580: dout <= { 2'd1, 8'd058, 10'd014 }; 
        'd1581: dout <= { 2'd1, 8'd037, 10'd208 }; 
        'd1582: dout <= { 2'd1, 8'd017, 10'd352 }; 
        'd1583: dout <= { 2'd2, 8'd059, 10'd197 }; 
        'd1584: dout <= { 2'd1, 8'd002, 10'd257 }; 
        'd1585: dout <= { 2'd1, 8'd060, 10'd308 }; 
        'd1586: dout <= { 2'd1, 8'd032, 10'd290 }; 
        'd1587: dout <= { 2'd1, 8'd024, 10'd124 }; 
        'd1588: dout <= { 2'd1, 8'd021, 10'd075 }; 
        'd1589: dout <= { 2'd1, 8'd067, 10'd217 }; 
        'd1590: dout <= { 2'd1, 8'd006, 10'd085 }; 
        'd1591: dout <= { 2'd1, 8'd067, 10'd299 }; 
        'd1592: dout <= { 2'd1, 8'd068, 10'd006 }; 
        'd1593: dout <= { 2'd1, 8'd064, 10'd095 }; 
        'd1594: dout <= { 2'd1, 8'd027, 10'd181 }; 
        'd1595: dout <= { 2'd2, 8'd034, 10'd094 }; 
        'd1596: dout <= { 2'd1, 8'd009, 10'd117 }; 
        'd1597: dout <= { 2'd1, 8'd014, 10'd065 }; 
        'd1598: dout <= { 2'd1, 8'd052, 10'd076 }; 
        'd1599: dout <= { 2'd1, 8'd032, 10'd197 }; 
        'd1600: dout <= { 2'd1, 8'd013, 10'd051 }; 
        'd1601: dout <= { 2'd1, 8'd065, 10'd273 }; 
        'd1602: dout <= { 2'd1, 8'd004, 10'd353 }; 
        'd1603: dout <= { 2'd1, 8'd001, 10'd138 }; 
        'd1604: dout <= { 2'd1, 8'd053, 10'd330 }; 
        'd1605: dout <= { 2'd1, 8'd047, 10'd125 }; 
        'd1606: dout <= { 2'd1, 8'd019, 10'd356 }; 
        'd1607: dout <= { 2'd2, 8'd050, 10'd233 }; 
        'd1608: dout <= { 2'd1, 8'd044, 10'd298 }; 
        'd1609: dout <= { 2'd1, 8'd046, 10'd344 }; 
        'd1610: dout <= { 2'd1, 8'd008, 10'd088 }; 
        'd1611: dout <= { 2'd1, 8'd030, 10'd241 }; 
        'd1612: dout <= { 2'd1, 8'd008, 10'd098 }; 
        'd1613: dout <= { 2'd1, 8'd033, 10'd193 }; 
        'd1614: dout <= { 2'd1, 8'd044, 10'd055 }; 
        'd1615: dout <= { 2'd1, 8'd064, 10'd229 }; 
        'd1616: dout <= { 2'd1, 8'd002, 10'd178 }; 
        'd1617: dout <= { 2'd1, 8'd008, 10'd121 }; 
        'd1618: dout <= { 2'd1, 8'd030, 10'd073 }; 
        'd1619: dout <= { 2'd2, 8'd046, 10'd030 }; 
        'd1620: dout <= { 2'd1, 8'd053, 10'd312 }; 
        'd1621: dout <= { 2'd1, 8'd053, 10'd033 }; 
        'd1622: dout <= { 2'd1, 8'd057, 10'd264 }; 
        'd1623: dout <= { 2'd1, 8'd041, 10'd040 }; 
        'd1624: dout <= { 2'd1, 8'd011, 10'd300 }; 
        'd1625: dout <= { 2'd1, 8'd001, 10'd026 }; 
        'd1626: dout <= { 2'd1, 8'd019, 10'd104 }; 
        'd1627: dout <= { 2'd1, 8'd045, 10'd078 }; 
        'd1628: dout <= { 2'd1, 8'd038, 10'd319 }; 
        'd1629: dout <= { 2'd1, 8'd016, 10'd321 }; 
        'd1630: dout <= { 2'd1, 8'd023, 10'd285 }; 
        'd1631: dout <= { 2'd2, 8'd049, 10'd274 }; 
        'd1632: dout <= { 2'd1, 8'd042, 10'd024 }; 
        'd1633: dout <= { 2'd1, 8'd028, 10'd064 }; 
        'd1634: dout <= { 2'd1, 8'd020, 10'd290 }; 
        'd1635: dout <= { 2'd1, 8'd027, 10'd207 }; 
        'd1636: dout <= { 2'd1, 8'd031, 10'd128 }; 
        'd1637: dout <= { 2'd1, 8'd028, 10'd171 }; 
        'd1638: dout <= { 2'd1, 8'd064, 10'd152 }; 
        'd1639: dout <= { 2'd1, 8'd006, 10'd180 }; 
        'd1640: dout <= { 2'd1, 8'd007, 10'd062 }; 
        'd1641: dout <= { 2'd1, 8'd067, 10'd037 }; 
        'd1642: dout <= { 2'd1, 8'd029, 10'd228 }; 
        'd1643: dout <= { 2'd2, 8'd071, 10'd010 }; 
        'd1644: dout <= { 2'd1, 8'd011, 10'd092 }; 
        'd1645: dout <= { 2'd1, 8'd012, 10'd202 }; 
        'd1646: dout <= { 2'd1, 8'd001, 10'd262 }; 
        'd1647: dout <= { 2'd1, 8'd029, 10'd311 }; 
        'd1648: dout <= { 2'd1, 8'd020, 10'd307 }; 
        'd1649: dout <= { 2'd1, 8'd025, 10'd176 }; 
        'd1650: dout <= { 2'd1, 8'd011, 10'd136 }; 
        'd1651: dout <= { 2'd1, 8'd069, 10'd353 }; 
        'd1652: dout <= { 2'd1, 8'd040, 10'd107 }; 
        'd1653: dout <= { 2'd1, 8'd038, 10'd253 }; 
        'd1654: dout <= { 2'd1, 8'd009, 10'd157 }; 
        'd1655: dout <= { 2'd2, 8'd004, 10'd125 }; 
        'd1656: dout <= { 2'd1, 8'd038, 10'd277 }; 
        'd1657: dout <= { 2'd1, 8'd059, 10'd332 }; 
        'd1658: dout <= { 2'd1, 8'd048, 10'd262 }; 
        'd1659: dout <= { 2'd1, 8'd006, 10'd100 }; 
        'd1660: dout <= { 2'd1, 8'd044, 10'd173 }; 
        'd1661: dout <= { 2'd1, 8'd062, 10'd060 }; 
        'd1662: dout <= { 2'd1, 8'd051, 10'd278 }; 
        'd1663: dout <= { 2'd1, 8'd057, 10'd085 }; 
        'd1664: dout <= { 2'd1, 8'd055, 10'd291 }; 
        'd1665: dout <= { 2'd1, 8'd043, 10'd016 }; 
        'd1666: dout <= { 2'd1, 8'd003, 10'd327 }; 
        'd1667: dout <= { 2'd2, 8'd069, 10'd344 }; 
        'd1668: dout <= { 2'd1, 8'd036, 10'd010 }; 
        'd1669: dout <= { 2'd1, 8'd070, 10'd154 }; 
        'd1670: dout <= { 2'd1, 8'd030, 10'd203 }; 
        'd1671: dout <= { 2'd1, 8'd014, 10'd285 }; 
        'd1672: dout <= { 2'd1, 8'd047, 10'd050 }; 
        'd1673: dout <= { 2'd1, 8'd016, 10'd246 }; 
        'd1674: dout <= { 2'd1, 8'd012, 10'd162 }; 
        'd1675: dout <= { 2'd1, 8'd035, 10'd164 }; 
        'd1676: dout <= { 2'd1, 8'd049, 10'd179 }; 
        'd1677: dout <= { 2'd1, 8'd010, 10'd061 }; 
        'd1678: dout <= { 2'd1, 8'd053, 10'd114 }; 
        'd1679: dout <= { 2'd2, 8'd048, 10'd318 }; 
        'd1680: dout <= { 2'd1, 8'd018, 10'd129 }; 
        'd1681: dout <= { 2'd1, 8'd033, 10'd333 }; 
        'd1682: dout <= { 2'd1, 8'd004, 10'd139 }; 
        'd1683: dout <= { 2'd1, 8'd065, 10'd153 }; 
        'd1684: dout <= { 2'd1, 8'd002, 10'd052 }; 
        'd1685: dout <= { 2'd1, 8'd061, 10'd337 }; 
        'd1686: dout <= { 2'd1, 8'd068, 10'd111 }; 
        'd1687: dout <= { 2'd1, 8'd026, 10'd275 }; 
        'd1688: dout <= { 2'd1, 8'd050, 10'd011 }; 
        'd1689: dout <= { 2'd1, 8'd052, 10'd122 }; 
        'd1690: dout <= { 2'd1, 8'd018, 10'd040 }; 
        'd1691: dout <= { 2'd2, 8'd051, 10'd069 }; 
        'd1692: dout <= { 2'd1, 8'd015, 10'd105 }; 
        'd1693: dout <= { 2'd1, 8'd039, 10'd103 }; 
        'd1694: dout <= { 2'd1, 8'd044, 10'd350 }; 
        'd1695: dout <= { 2'd1, 8'd056, 10'd065 }; 
        'd1696: dout <= { 2'd1, 8'd000, 10'd200 }; 
        'd1697: dout <= { 2'd1, 8'd013, 10'd319 }; 
        'd1698: dout <= { 2'd1, 8'd071, 10'd076 }; 
        'd1699: dout <= { 2'd1, 8'd014, 10'd111 }; 
        'd1700: dout <= { 2'd1, 8'd011, 10'd336 }; 
        'd1701: dout <= { 2'd1, 8'd021, 10'd181 }; 
        'd1702: dout <= { 2'd1, 8'd040, 10'd015 }; 
        'd1703: dout <= { 2'd2, 8'd016, 10'd071 }; 
        'd1704: dout <= { 2'd1, 8'd026, 10'd048 }; 
        'd1705: dout <= { 2'd1, 8'd054, 10'd128 }; 
        'd1706: dout <= { 2'd1, 8'd027, 10'd181 }; 
        'd1707: dout <= { 2'd1, 8'd057, 10'd219 }; 
        'd1708: dout <= { 2'd1, 8'd037, 10'd103 }; 
        'd1709: dout <= { 2'd1, 8'd059, 10'd329 }; 
        'd1710: dout <= { 2'd1, 8'd056, 10'd050 }; 
        'd1711: dout <= { 2'd1, 8'd033, 10'd341 }; 
        'd1712: dout <= { 2'd1, 8'd054, 10'd229 }; 
        'd1713: dout <= { 2'd1, 8'd011, 10'd243 }; 
        'd1714: dout <= { 2'd1, 8'd070, 10'd311 }; 
        'd1715: dout <= { 2'd2, 8'd054, 10'd203 }; 
        'd1716: dout <= { 2'd1, 8'd003, 10'd217 }; 
        'd1717: dout <= { 2'd1, 8'd026, 10'd212 }; 
        'd1718: dout <= { 2'd1, 8'd022, 10'd058 }; 
        'd1719: dout <= { 2'd1, 8'd068, 10'd315 }; 
        'd1720: dout <= { 2'd1, 8'd010, 10'd081 }; 
        'd1721: dout <= { 2'd1, 8'd003, 10'd186 }; 
        'd1722: dout <= { 2'd1, 8'd014, 10'd332 }; 
        'd1723: dout <= { 2'd1, 8'd065, 10'd235 }; 
        'd1724: dout <= { 2'd1, 8'd025, 10'd207 }; 
        'd1725: dout <= { 2'd1, 8'd054, 10'd051 }; 
        'd1726: dout <= { 2'd1, 8'd006, 10'd352 }; 
        'd1727: dout <= { 2'd2, 8'd037, 10'd335 }; 
        'd1728: dout <= { 2'd1, 8'd056, 10'd345 }; 
        'd1729: dout <= { 2'd1, 8'd021, 10'd227 }; 
        'd1730: dout <= { 2'd1, 8'd007, 10'd228 }; 
        'd1731: dout <= { 2'd1, 8'd069, 10'd186 }; 
        'd1732: dout <= { 2'd1, 8'd055, 10'd230 }; 
        'd1733: dout <= { 2'd1, 8'd043, 10'd112 }; 
        'd1734: dout <= { 2'd1, 8'd045, 10'd343 }; 
        'd1735: dout <= { 2'd1, 8'd004, 10'd050 }; 
        'd1736: dout <= { 2'd1, 8'd056, 10'd359 }; 
        'd1737: dout <= { 2'd1, 8'd004, 10'd121 }; 
        'd1738: dout <= { 2'd1, 8'd028, 10'd133 }; 
        'd1739: dout <= { 2'd2, 8'd061, 10'd282 }; 
        'd1740: dout <= { 2'd1, 8'd057, 10'd051 }; 
        'd1741: dout <= { 2'd1, 8'd037, 10'd239 }; 
        'd1742: dout <= { 2'd1, 8'd016, 10'd256 }; 
        'd1743: dout <= { 2'd1, 8'd070, 10'd136 }; 
        'd1744: dout <= { 2'd1, 8'd023, 10'd289 }; 
        'd1745: dout <= { 2'd1, 8'd054, 10'd351 }; 
        'd1746: dout <= { 2'd1, 8'd069, 10'd284 }; 
        'd1747: dout <= { 2'd1, 8'd066, 10'd341 }; 
        'd1748: dout <= { 2'd1, 8'd034, 10'd184 }; 
        'd1749: dout <= { 2'd1, 8'd059, 10'd070 }; 
        'd1750: dout <= { 2'd1, 8'd071, 10'd196 }; 
        'd1751: dout <= { 2'd2, 8'd020, 10'd122 }; 
        'd1752: dout <= { 2'd1, 8'd039, 10'd228 }; 
        'd1753: dout <= { 2'd1, 8'd006, 10'd245 }; 
        'd1754: dout <= { 2'd1, 8'd040, 10'd213 }; 
        'd1755: dout <= { 2'd1, 8'd050, 10'd252 }; 
        'd1756: dout <= { 2'd1, 8'd040, 10'd354 }; 
        'd1757: dout <= { 2'd1, 8'd049, 10'd024 }; 
        'd1758: dout <= { 2'd1, 8'd018, 10'd084 }; 
        'd1759: dout <= { 2'd1, 8'd039, 10'd303 }; 
        'd1760: dout <= { 2'd1, 8'd044, 10'd199 }; 
        'd1761: dout <= { 2'd1, 8'd061, 10'd173 }; 
        'd1762: dout <= { 2'd1, 8'd024, 10'd062 }; 
        'd1763: dout <= { 2'd2, 8'd066, 10'd242 }; 
        'd1764: dout <= { 2'd1, 8'd032, 10'd019 }; 
        'd1765: dout <= { 2'd1, 8'd071, 10'd112 }; 
        'd1766: dout <= { 2'd1, 8'd047, 10'd324 }; 
        'd1767: dout <= { 2'd1, 8'd071, 10'd289 }; 
        'd1768: dout <= { 2'd1, 8'd052, 10'd117 }; 
        'd1769: dout <= { 2'd1, 8'd052, 10'd056 }; 
        'd1770: dout <= { 2'd1, 8'd048, 10'd179 }; 
        'd1771: dout <= { 2'd1, 8'd048, 10'd354 }; 
        'd1772: dout <= { 2'd1, 8'd061, 10'd309 }; 
        'd1773: dout <= { 2'd1, 8'd022, 10'd230 }; 
        'd1774: dout <= { 2'd1, 8'd066, 10'd088 }; 
        'd1775: dout <= { 2'd2, 8'd024, 10'd338 }; 
        'd1776: dout <= { 2'd1, 8'd063, 10'd348 }; 
        'd1777: dout <= { 2'd1, 8'd042, 10'd327 }; 
        'd1778: dout <= { 2'd1, 8'd056, 10'd001 }; 
        'd1779: dout <= { 2'd1, 8'd009, 10'd066 }; 
        'd1780: dout <= { 2'd1, 8'd003, 10'd145 }; 
        'd1781: dout <= { 2'd1, 8'd000, 10'd313 }; 
        'd1782: dout <= { 2'd1, 8'd039, 10'd119 }; 
        'd1783: dout <= { 2'd1, 8'd032, 10'd135 }; 
        'd1784: dout <= { 2'd1, 8'd030, 10'd353 }; 
        'd1785: dout <= { 2'd1, 8'd005, 10'd209 }; 
        'd1786: dout <= { 2'd1, 8'd056, 10'd025 }; 
        'd1787: dout <= { 2'd2, 8'd008, 10'd056 }; 
        'd1788: dout <= { 2'd1, 8'd017, 10'd005 }; 
        'd1789: dout <= { 2'd1, 8'd064, 10'd293 }; 
        'd1790: dout <= { 2'd1, 8'd010, 10'd187 }; 
        'd1791: dout <= { 2'd1, 8'd051, 10'd075 }; 
        'd1792: dout <= { 2'd1, 8'd034, 10'd238 }; 
        'd1793: dout <= { 2'd1, 8'd034, 10'd082 }; 
        'd1794: dout <= { 2'd1, 8'd032, 10'd142 }; 
        'd1795: dout <= { 2'd1, 8'd020, 10'd166 }; 
        'd1796: dout <= { 2'd1, 8'd018, 10'd336 }; 
        'd1797: dout <= { 2'd1, 8'd049, 10'd247 }; 
        'd1798: dout <= { 2'd1, 8'd015, 10'd306 }; 
        'd1799: dout <= { 2'd2, 8'd052, 10'd223 }; 
        'd1800: dout <= { 2'd1, 8'd043, 10'd181 }; 
        'd1801: dout <= { 2'd1, 8'd000, 10'd134 }; 
        'd1802: dout <= { 2'd1, 8'd066, 10'd340 }; 
        'd1803: dout <= { 2'd1, 8'd046, 10'd182 }; 
        'd1804: dout <= { 2'd1, 8'd035, 10'd331 }; 
        'd1805: dout <= { 2'd1, 8'd037, 10'd101 }; 
        'd1806: dout <= { 2'd1, 8'd070, 10'd274 }; 
        'd1807: dout <= { 2'd1, 8'd036, 10'd041 }; 
        'd1808: dout <= { 2'd1, 8'd010, 10'd234 }; 
        'd1809: dout <= { 2'd1, 8'd001, 10'd067 }; 
        'd1810: dout <= { 2'd1, 8'd046, 10'd332 }; 
        'd1811: dout <= { 2'd2, 8'd005, 10'd210 }; 
        'd1812: dout <= { 2'd1, 8'd006, 10'd285 }; 
        'd1813: dout <= { 2'd1, 8'd025, 10'd049 }; 
        'd1814: dout <= { 2'd1, 8'd005, 10'd160 }; 
        'd1815: dout <= { 2'd1, 8'd038, 10'd324 }; 
        'd1816: dout <= { 2'd1, 8'd004, 10'd034 }; 
        'd1817: dout <= { 2'd1, 8'd058, 10'd244 }; 
        'd1818: dout <= { 2'd1, 8'd041, 10'd267 }; 
        'd1819: dout <= { 2'd1, 8'd012, 10'd280 }; 
        'd1820: dout <= { 2'd1, 8'd060, 10'd250 }; 
        'd1821: dout <= { 2'd1, 8'd041, 10'd341 }; 
        'd1822: dout <= { 2'd1, 8'd007, 10'd184 }; 
        'd1823: dout <= { 2'd2, 8'd040, 10'd021 }; 
        'd1824: dout <= { 2'd1, 8'd047, 10'd261 }; 
        'd1825: dout <= { 2'd1, 8'd036, 10'd293 }; 
        'd1826: dout <= { 2'd1, 8'd031, 10'd279 }; 
        'd1827: dout <= { 2'd1, 8'd022, 10'd211 }; 
        'd1828: dout <= { 2'd1, 8'd017, 10'd204 }; 
        'd1829: dout <= { 2'd1, 8'd040, 10'd098 }; 
        'd1830: dout <= { 2'd1, 8'd022, 10'd141 }; 
        'd1831: dout <= { 2'd1, 8'd047, 10'd078 }; 
        'd1832: dout <= { 2'd1, 8'd003, 10'd259 }; 
        'd1833: dout <= { 2'd1, 8'd044, 10'd273 }; 
        'd1834: dout <= { 2'd1, 8'd068, 10'd173 }; 
        'd1835: dout <= { 2'd2, 8'd065, 10'd194 }; 
        'd1836: dout <= { 2'd1, 8'd023, 10'd057 }; 
        'd1837: dout <= { 2'd1, 8'd019, 10'd041 }; 
        'd1838: dout <= { 2'd1, 8'd003, 10'd243 }; 
        'd1839: dout <= { 2'd1, 8'd015, 10'd226 }; 
        'd1840: dout <= { 2'd1, 8'd048, 10'd310 }; 
        'd1841: dout <= { 2'd1, 8'd007, 10'd298 }; 
        'd1842: dout <= { 2'd1, 8'd023, 10'd110 }; 
        'd1843: dout <= { 2'd1, 8'd016, 10'd262 }; 
        'd1844: dout <= { 2'd1, 8'd023, 10'd077 }; 
        'd1845: dout <= { 2'd1, 8'd055, 10'd111 }; 
        'd1846: dout <= { 2'd1, 8'd035, 10'd324 }; 
        'd1847: dout <= { 2'd2, 8'd029, 10'd094 }; 
        'd1848: dout <= { 2'd1, 8'd067, 10'd147 }; 
        'd1849: dout <= { 2'd1, 8'd063, 10'd339 }; 
        'd1850: dout <= { 2'd1, 8'd069, 10'd198 }; 
        'd1851: dout <= { 2'd1, 8'd049, 10'd056 }; 
        'd1852: dout <= { 2'd1, 8'd058, 10'd100 }; 
        'd1853: dout <= { 2'd1, 8'd053, 10'd068 }; 
        'd1854: dout <= { 2'd1, 8'd060, 10'd097 }; 
        'd1855: dout <= { 2'd1, 8'd070, 10'd014 }; 
        'd1856: dout <= { 2'd1, 8'd005, 10'd011 }; 
        'd1857: dout <= { 2'd1, 8'd014, 10'd318 }; 
        'd1858: dout <= { 2'd1, 8'd026, 10'd284 }; 
        'd1859: dout <= { 2'd2, 8'd070, 10'd059 }; 
        'd1860: dout <= { 2'd1, 8'd062, 10'd296 }; 
        'd1861: dout <= { 2'd1, 8'd055, 10'd183 }; 
        'd1862: dout <= { 2'd1, 8'd017, 10'd319 }; 
        'd1863: dout <= { 2'd1, 8'd016, 10'd070 }; 
        'd1864: dout <= { 2'd1, 8'd005, 10'd053 }; 
        'd1865: dout <= { 2'd1, 8'd030, 10'd329 }; 
        'd1866: dout <= { 2'd1, 8'd066, 10'd196 }; 
        'd1867: dout <= { 2'd1, 8'd042, 10'd138 }; 
        'd1868: dout <= { 2'd1, 8'd022, 10'd264 }; 
        'd1869: dout <= { 2'd1, 8'd050, 10'd327 }; 
        'd1870: dout <= { 2'd1, 8'd039, 10'd123 }; 
        'd1871: dout <= { 2'd2, 8'd014, 10'd352 }; 
        'd1872: dout <= { 2'd1, 8'd007, 10'd086 }; 
        'd1873: dout <= { 2'd1, 8'd024, 10'd306 }; 
        'd1874: dout <= { 2'd1, 8'd045, 10'd107 }; 
        'd1875: dout <= { 2'd1, 8'd062, 10'd184 }; 
        'd1876: dout <= { 2'd1, 8'd039, 10'd055 }; 
        'd1877: dout <= { 2'd1, 8'd009, 10'd329 }; 
        'd1878: dout <= { 2'd1, 8'd029, 10'd228 }; 
        'd1879: dout <= { 2'd1, 8'd028, 10'd314 }; 
        'd1880: dout <= { 2'd1, 8'd041, 10'd072 }; 
        'd1881: dout <= { 2'd1, 8'd045, 10'd311 }; 
        'd1882: dout <= { 2'd1, 8'd033, 10'd335 }; 
        'd1883: dout <= { 2'd2, 8'd010, 10'd131 }; 
        'd1884: dout <= { 2'd1, 8'd058, 10'd110 }; 
        'd1885: dout <= { 2'd1, 8'd009, 10'd169 }; 
        'd1886: dout <= { 2'd1, 8'd013, 10'd040 }; 
        'd1887: dout <= { 2'd1, 8'd042, 10'd288 }; 
        'd1888: dout <= { 2'd1, 8'd007, 10'd044 }; 
        'd1889: dout <= { 2'd1, 8'd005, 10'd120 }; 
        'd1890: dout <= { 2'd1, 8'd055, 10'd164 }; 
        'd1891: dout <= { 2'd1, 8'd071, 10'd341 }; 
        'd1892: dout <= { 2'd1, 8'd015, 10'd143 }; 
        'd1893: dout <= { 2'd1, 8'd063, 10'd357 }; 
        'd1894: dout <= { 2'd1, 8'd065, 10'd236 }; 
        'd1895: dout <= { 2'd2, 8'd019, 10'd051 }; 
        'd1896: dout <= { 2'd1, 8'd025, 10'd284 }; 
        'd1897: dout <= { 2'd1, 8'd062, 10'd156 }; 
        'd1898: dout <= { 2'd1, 8'd050, 10'd137 }; 
        'd1899: dout <= { 2'd1, 8'd063, 10'd316 }; 
        'd1900: dout <= { 2'd1, 8'd054, 10'd035 }; 
        'd1901: dout <= { 2'd1, 8'd015, 10'd117 }; 
        'd1902: dout <= { 2'd1, 8'd027, 10'd051 }; 
        'd1903: dout <= { 2'd1, 8'd031, 10'd075 }; 
        'd1904: dout <= { 2'd1, 8'd000, 10'd345 }; 
        'd1905: dout <= { 2'd1, 8'd020, 10'd304 }; 
        'd1906: dout <= { 2'd1, 8'd032, 10'd223 }; 
        'd1907: dout <= { 2'd2, 8'd028, 10'd253 }; 
        'd1908: dout <= { 2'd1, 8'd000, 10'd114 }; 
        'd1909: dout <= { 2'd1, 8'd067, 10'd079 }; 
        'd1910: dout <= { 2'd1, 8'd051, 10'd264 }; 
        'd1911: dout <= { 2'd1, 8'd045, 10'd118 }; 
        'd1912: dout <= { 2'd1, 8'd012, 10'd346 }; 
        'd1913: dout <= { 2'd1, 8'd046, 10'd089 }; 
        'd1914: dout <= { 2'd1, 8'd002, 10'd156 }; 
        'd1915: dout <= { 2'd1, 8'd052, 10'd145 }; 
        'd1916: dout <= { 2'd1, 8'd062, 10'd227 }; 
        'd1917: dout <= { 2'd1, 8'd031, 10'd150 }; 
        'd1918: dout <= { 2'd1, 8'd060, 10'd158 }; 
        'd1919: dout <= { 2'd2, 8'd001, 10'd134 }; 
        'd1920: dout <= { 2'd1, 8'd064, 10'd225 }; 
        'd1921: dout <= { 2'd1, 8'd043, 10'd156 }; 
        'd1922: dout <= { 2'd1, 8'd041, 10'd346 }; 
        'd1923: dout <= { 2'd1, 8'd043, 10'd032 }; 
        'd1924: dout <= { 2'd1, 8'd067, 10'd175 }; 
        'd1925: dout <= { 2'd1, 8'd038, 10'd266 }; 
        'd1926: dout <= { 2'd1, 8'd057, 10'd100 }; 
        'd1927: dout <= { 2'd1, 8'd046, 10'd099 }; 
        'd1928: dout <= { 2'd1, 8'd051, 10'd344 }; 
        'd1929: dout <= { 2'd1, 8'd058, 10'd040 }; 
        'd1930: dout <= { 2'd1, 8'd002, 10'd035 }; 
        'd1931: dout <= { 2'd2, 8'd013, 10'd163 }; 
        'd1932: dout <= { 2'd1, 8'd028, 10'd050 }; 
        'd1933: dout <= { 2'd1, 8'd065, 10'd082 }; 
        'd1934: dout <= { 2'd1, 8'd038, 10'd192 }; 
        'd1935: dout <= { 2'd1, 8'd026, 10'd021 }; 
        'd1936: dout <= { 2'd1, 8'd064, 10'd321 }; 
        'd1937: dout <= { 2'd1, 8'd017, 10'd088 }; 
        'd1938: dout <= { 2'd1, 8'd047, 10'd039 }; 
        'd1939: dout <= { 2'd1, 8'd008, 10'd246 }; 
        'd1940: dout <= { 2'd1, 8'd024, 10'd034 }; 
        'd1941: dout <= { 2'd1, 8'd012, 10'd103 }; 
        'd1942: dout <= { 2'd1, 8'd069, 10'd007 }; 
        'd1943: dout <= { 2'd2, 8'd060, 10'd208 }; 
        'd1944: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd1945: dout <= { 2'd1, 8'd035, 10'd257 }; 
        'd1946: dout <= { 2'd2, 8'd013, 10'd259 }; 
        'd1947: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd1948: dout <= { 2'd1, 8'd062, 10'd145 }; 
        'd1949: dout <= { 2'd2, 8'd050, 10'd041 }; 
        'd1950: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd1951: dout <= { 2'd1, 8'd008, 10'd130 }; 
        'd1952: dout <= { 2'd2, 8'd033, 10'd149 }; 
        'd1953: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd1954: dout <= { 2'd1, 8'd059, 10'd170 }; 
        'd1955: dout <= { 2'd2, 8'd052, 10'd108 }; 
        'd1956: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd1957: dout <= { 2'd1, 8'd000, 10'd209 }; 
        'd1958: dout <= { 2'd2, 8'd042, 10'd185 }; 
        'd1959: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd1960: dout <= { 2'd1, 8'd012, 10'd256 }; 
        'd1961: dout <= { 2'd2, 8'd016, 10'd342 }; 
        'd1962: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd1963: dout <= { 2'd1, 8'd039, 10'd288 }; 
        'd1964: dout <= { 2'd2, 8'd023, 10'd266 }; 
        'd1965: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd1966: dout <= { 2'd1, 8'd034, 10'd263 }; 
        'd1967: dout <= { 2'd2, 8'd027, 10'd152 }; 
        'd1968: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd1969: dout <= { 2'd1, 8'd001, 10'd074 }; 
        'd1970: dout <= { 2'd2, 8'd038, 10'd277 }; 
        'd1971: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd1972: dout <= { 2'd1, 8'd064, 10'd156 }; 
        'd1973: dout <= { 2'd2, 8'd007, 10'd259 }; 
        'd1974: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd1975: dout <= { 2'd1, 8'd070, 10'd208 }; 
        'd1976: dout <= { 2'd2, 8'd067, 10'd286 }; 
        'd1977: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd1978: dout <= { 2'd1, 8'd028, 10'd101 }; 
        'd1979: dout <= { 2'd2, 8'd036, 10'd307 }; 
        'd1980: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd1981: dout <= { 2'd1, 8'd069, 10'd305 }; 
        'd1982: dout <= { 2'd2, 8'd005, 10'd201 }; 
        'd1983: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd1984: dout <= { 2'd1, 8'd041, 10'd154 }; 
        'd1985: dout <= { 2'd2, 8'd022, 10'd010 }; 
        'd1986: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd1987: dout <= { 2'd1, 8'd006, 10'd184 }; 
        'd1988: dout <= { 2'd2, 8'd061, 10'd191 }; 
        'd1989: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd1990: dout <= { 2'd1, 8'd010, 10'd267 }; 
        'd1991: dout <= { 2'd2, 8'd025, 10'd184 }; 
        'd1992: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd1993: dout <= { 2'd1, 8'd031, 10'd084 }; 
        'd1994: dout <= { 2'd2, 8'd026, 10'd293 }; 
        'd1995: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd1996: dout <= { 2'd1, 8'd030, 10'd316 }; 
        'd1997: dout <= { 2'd2, 8'd068, 10'd080 }; 
        'd1998: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd1999: dout <= { 2'd1, 8'd047, 10'd274 }; 
        'd2000: dout <= { 2'd2, 8'd071, 10'd058 }; 
        'd2001: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd2002: dout <= { 2'd1, 8'd004, 10'd023 }; 
        'd2003: dout <= { 2'd2, 8'd045, 10'd269 }; 
        'd2004: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd2005: dout <= { 2'd1, 8'd011, 10'd061 }; 
        'd2006: dout <= { 2'd2, 8'd049, 10'd050 }; 
        'd2007: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd2008: dout <= { 2'd1, 8'd051, 10'd185 }; 
        'd2009: dout <= { 2'd2, 8'd003, 10'd359 }; 
        'd2010: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd2011: dout <= { 2'd1, 8'd018, 10'd316 }; 
        'd2012: dout <= { 2'd2, 8'd040, 10'd302 }; 
        'd2013: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd2014: dout <= { 2'd1, 8'd029, 10'd149 }; 
        'd2015: dout <= { 2'd2, 8'd019, 10'd196 }; 
        'd2016: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd2017: dout <= { 2'd1, 8'd015, 10'd223 }; 
        'd2018: dout <= { 2'd2, 8'd017, 10'd300 }; 
        'd2019: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd2020: dout <= { 2'd1, 8'd057, 10'd088 }; 
        'd2021: dout <= { 2'd2, 8'd053, 10'd051 }; 
        'd2022: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd2023: dout <= { 2'd1, 8'd021, 10'd008 }; 
        'd2024: dout <= { 2'd2, 8'd024, 10'd277 }; 
        'd2025: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd2026: dout <= { 2'd1, 8'd055, 10'd079 }; 
        'd2027: dout <= { 2'd2, 8'd020, 10'd112 }; 
        'd2028: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd2029: dout <= { 2'd1, 8'd002, 10'd094 }; 
        'd2030: dout <= { 2'd2, 8'd044, 10'd132 }; 
        'd2031: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd2032: dout <= { 2'd1, 8'd037, 10'd059 }; 
        'd2033: dout <= { 2'd2, 8'd046, 10'd243 }; 
        'd2034: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd2035: dout <= { 2'd1, 8'd032, 10'd188 }; 
        'd2036: dout <= { 2'd2, 8'd063, 10'd313 }; 
        'd2037: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd2038: dout <= { 2'd1, 8'd058, 10'd024 }; 
        'd2039: dout <= { 2'd2, 8'd009, 10'd064 }; 
        'd2040: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd2041: dout <= { 2'd1, 8'd054, 10'd322 }; 
        'd2042: dout <= { 2'd2, 8'd056, 10'd161 }; 
        'd2043: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd2044: dout <= { 2'd1, 8'd043, 10'd272 }; 
        'd2045: dout <= { 2'd2, 8'd014, 10'd028 }; 
        'd2046: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd2047: dout <= { 2'd1, 8'd065, 10'd188 }; 
        'd2048: dout <= { 2'd2, 8'd066, 10'd186 }; 
        'd2049: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd2050: dout <= { 2'd1, 8'd060, 10'd190 }; 
        'd2051: dout <= { 2'd2, 8'd048, 10'd240 }; 
        'd2052: dout <= { 2'd1, 8'd036, 10'd000 }; 
        'd2053: dout <= { 2'd1, 8'd028, 10'd347 }; 
        'd2054: dout <= { 2'd2, 8'd048, 10'd193 }; 
        'd2055: dout <= { 2'd1, 8'd037, 10'd000 }; 
        'd2056: dout <= { 2'd1, 8'd049, 10'd312 }; 
        'd2057: dout <= { 2'd2, 8'd063, 10'd092 }; 
        'd2058: dout <= { 2'd1, 8'd038, 10'd000 }; 
        'd2059: dout <= { 2'd1, 8'd038, 10'd068 }; 
        'd2060: dout <= { 2'd2, 8'd059, 10'd174 }; 
        'd2061: dout <= { 2'd1, 8'd039, 10'd000 }; 
        'd2062: dout <= { 2'd1, 8'd029, 10'd294 }; 
        'd2063: dout <= { 2'd2, 8'd021, 10'd071 }; 
        'd2064: dout <= { 2'd1, 8'd040, 10'd000 }; 
        'd2065: dout <= { 2'd1, 8'd025, 10'd315 }; 
        'd2066: dout <= { 2'd2, 8'd026, 10'd096 }; 
        'd2067: dout <= { 2'd1, 8'd041, 10'd000 }; 
        'd2068: dout <= { 2'd1, 8'd046, 10'd104 }; 
        'd2069: dout <= { 2'd2, 8'd009, 10'd342 }; 
        'd2070: dout <= { 2'd1, 8'd042, 10'd000 }; 
        'd2071: dout <= { 2'd1, 8'd064, 10'd338 }; 
        'd2072: dout <= { 2'd2, 8'd053, 10'd177 }; 
        'd2073: dout <= { 2'd1, 8'd043, 10'd000 }; 
        'd2074: dout <= { 2'd1, 8'd023, 10'd304 }; 
        'd2075: dout <= { 2'd2, 8'd008, 10'd357 }; 
        'd2076: dout <= { 2'd1, 8'd044, 10'd000 }; 
        'd2077: dout <= { 2'd1, 8'd015, 10'd167 }; 
        'd2078: dout <= { 2'd2, 8'd060, 10'd015 }; 
        'd2079: dout <= { 2'd1, 8'd045, 10'd000 }; 
        'd2080: dout <= { 2'd1, 8'd042, 10'd337 }; 
        'd2081: dout <= { 2'd2, 8'd013, 10'd014 }; 
        'd2082: dout <= { 2'd1, 8'd046, 10'd000 }; 
        'd2083: dout <= { 2'd1, 8'd044, 10'd194 }; 
        'd2084: dout <= { 2'd2, 8'd011, 10'd288 }; 
        'd2085: dout <= { 2'd1, 8'd047, 10'd000 }; 
        'd2086: dout <= { 2'd1, 8'd033, 10'd156 }; 
        'd2087: dout <= { 2'd2, 8'd027, 10'd211 }; 
        'd2088: dout <= { 2'd1, 8'd048, 10'd000 }; 
        'd2089: dout <= { 2'd1, 8'd062, 10'd064 }; 
        'd2090: dout <= { 2'd2, 8'd051, 10'd215 }; 
        'd2091: dout <= { 2'd1, 8'd049, 10'd000 }; 
        'd2092: dout <= { 2'd1, 8'd057, 10'd130 }; 
        'd2093: dout <= { 2'd2, 8'd031, 10'd199 }; 
        'd2094: dout <= { 2'd1, 8'd050, 10'd000 }; 
        'd2095: dout <= { 2'd1, 8'd039, 10'd033 }; 
        'd2096: dout <= { 2'd2, 8'd024, 10'd090 }; 
        'd2097: dout <= { 2'd1, 8'd051, 10'd000 }; 
        'd2098: dout <= { 2'd1, 8'd052, 10'd346 }; 
        'd2099: dout <= { 2'd2, 8'd066, 10'd342 }; 
        'd2100: dout <= { 2'd1, 8'd052, 10'd000 }; 
        'd2101: dout <= { 2'd1, 8'd043, 10'd200 }; 
        'd2102: dout <= { 2'd2, 8'd032, 10'd122 }; 
        'd2103: dout <= { 2'd1, 8'd053, 10'd000 }; 
        'd2104: dout <= { 2'd1, 8'd014, 10'd096 }; 
        'd2105: dout <= { 2'd2, 8'd067, 10'd017 }; 
        'd2106: dout <= { 2'd1, 8'd054, 10'd000 }; 
        'd2107: dout <= { 2'd1, 8'd017, 10'd086 }; 
        'd2108: dout <= { 2'd2, 8'd070, 10'd288 }; 
        'd2109: dout <= { 2'd1, 8'd055, 10'd000 }; 
        'd2110: dout <= { 2'd1, 8'd019, 10'd193 }; 
        'd2111: dout <= { 2'd2, 8'd047, 10'd056 }; 
        'd2112: dout <= { 2'd1, 8'd056, 10'd000 }; 
        'd2113: dout <= { 2'd1, 8'd002, 10'd339 }; 
        'd2114: dout <= { 2'd2, 8'd020, 10'd183 }; 
        'd2115: dout <= { 2'd1, 8'd057, 10'd000 }; 
        'd2116: dout <= { 2'd1, 8'd041, 10'd187 }; 
        'd2117: dout <= { 2'd2, 8'd069, 10'd084 }; 
        'd2118: dout <= { 2'd1, 8'd058, 10'd000 }; 
        'd2119: dout <= { 2'd1, 8'd005, 10'd137 }; 
        'd2120: dout <= { 2'd2, 8'd012, 10'd114 }; 
        'd2121: dout <= { 2'd1, 8'd059, 10'd000 }; 
        'd2122: dout <= { 2'd1, 8'd058, 10'd021 }; 
        'd2123: dout <= { 2'd2, 8'd068, 10'd083 }; 
        'd2124: dout <= { 2'd1, 8'd060, 10'd000 }; 
        'd2125: dout <= { 2'd1, 8'd004, 10'd358 }; 
        'd2126: dout <= { 2'd2, 8'd035, 10'd241 }; 
        'd2127: dout <= { 2'd1, 8'd061, 10'd000 }; 
        'd2128: dout <= { 2'd1, 8'd007, 10'd287 }; 
        'd2129: dout <= { 2'd2, 8'd001, 10'd346 }; 
        'd2130: dout <= { 2'd1, 8'd062, 10'd000 }; 
        'd2131: dout <= { 2'd1, 8'd006, 10'd341 }; 
        'd2132: dout <= { 2'd2, 8'd071, 10'd285 }; 
        'd2133: dout <= { 2'd1, 8'd063, 10'd000 }; 
        'd2134: dout <= { 2'd1, 8'd018, 10'd172 }; 
        'd2135: dout <= { 2'd2, 8'd030, 10'd051 }; 
        'd2136: dout <= { 2'd1, 8'd064, 10'd000 }; 
        'd2137: dout <= { 2'd1, 8'd034, 10'd115 }; 
        'd2138: dout <= { 2'd2, 8'd061, 10'd018 }; 
        'd2139: dout <= { 2'd1, 8'd065, 10'd000 }; 
        'd2140: dout <= { 2'd1, 8'd055, 10'd278 }; 
        'd2141: dout <= { 2'd2, 8'd000, 10'd203 }; 
        'd2142: dout <= { 2'd1, 8'd066, 10'd000 }; 
        'd2143: dout <= { 2'd1, 8'd022, 10'd236 }; 
        'd2144: dout <= { 2'd2, 8'd016, 10'd051 }; 
        'd2145: dout <= { 2'd1, 8'd067, 10'd000 }; 
        'd2146: dout <= { 2'd1, 8'd037, 10'd275 }; 
        'd2147: dout <= { 2'd2, 8'd010, 10'd013 }; 
        'd2148: dout <= { 2'd1, 8'd068, 10'd000 }; 
        'd2149: dout <= { 2'd1, 8'd003, 10'd211 }; 
        'd2150: dout <= { 2'd2, 8'd040, 10'd168 }; 
        'd2151: dout <= { 2'd1, 8'd069, 10'd000 }; 
        'd2152: dout <= { 2'd1, 8'd054, 10'd107 }; 
        'd2153: dout <= { 2'd2, 8'd056, 10'd316 }; 
        'd2154: dout <= { 2'd1, 8'd070, 10'd000 }; 
        'd2155: dout <= { 2'd1, 8'd036, 10'd049 }; 
        'd2156: dout <= { 2'd2, 8'd045, 10'd040 }; 
        'd2157: dout <= { 2'd1, 8'd071, 10'd000 }; 
        'd2158: dout <= { 2'd1, 8'd050, 10'd047 }; 
        'd2159: dout <= { 2'd3, 8'd065, 10'd107 }; 
        // Q=60, BaseAddr=2160
        'd2160: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd2161: dout <= { 2'd1, 8'd051, 10'd174 }; 
        'd2162: dout <= { 2'd1, 8'd023, 10'd267 }; 
        'd2163: dout <= { 2'd1, 8'd026, 10'd008 }; 
        'd2164: dout <= { 2'd1, 8'd046, 10'd213 }; 
        'd2165: dout <= { 2'd1, 8'd025, 10'd134 }; 
        'd2166: dout <= { 2'd1, 8'd006, 10'd137 }; 
        'd2167: dout <= { 2'd1, 8'd007, 10'd046 }; 
        'd2168: dout <= { 2'd1, 8'd000, 10'd004 }; 
        'd2169: dout <= { 2'd1, 8'd013, 10'd311 }; 
        'd2170: dout <= { 2'd1, 8'd039, 10'd154 }; 
        'd2171: dout <= { 2'd1, 8'd019, 10'd176 }; 
        'd2172: dout <= { 2'd2, 8'd048, 10'd348 }; 
        'd2173: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd2174: dout <= { 2'd1, 8'd059, 10'd296 }; 
        'd2175: dout <= { 2'd1, 8'd033, 10'd138 }; 
        'd2176: dout <= { 2'd1, 8'd013, 10'd107 }; 
        'd2177: dout <= { 2'd1, 8'd044, 10'd103 }; 
        'd2178: dout <= { 2'd1, 8'd020, 10'd085 }; 
        'd2179: dout <= { 2'd1, 8'd004, 10'd097 }; 
        'd2180: dout <= { 2'd1, 8'd032, 10'd213 }; 
        'd2181: dout <= { 2'd1, 8'd027, 10'd286 }; 
        'd2182: dout <= { 2'd1, 8'd040, 10'd165 }; 
        'd2183: dout <= { 2'd1, 8'd007, 10'd224 }; 
        'd2184: dout <= { 2'd1, 8'd025, 10'd230 }; 
        'd2185: dout <= { 2'd2, 8'd003, 10'd308 }; 
        'd2186: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd2187: dout <= { 2'd1, 8'd017, 10'd299 }; 
        'd2188: dout <= { 2'd1, 8'd024, 10'd100 }; 
        'd2189: dout <= { 2'd1, 8'd041, 10'd144 }; 
        'd2190: dout <= { 2'd1, 8'd028, 10'd310 }; 
        'd2191: dout <= { 2'd1, 8'd014, 10'd213 }; 
        'd2192: dout <= { 2'd1, 8'd035, 10'd098 }; 
        'd2193: dout <= { 2'd1, 8'd056, 10'd242 }; 
        'd2194: dout <= { 2'd1, 8'd050, 10'd182 }; 
        'd2195: dout <= { 2'd1, 8'd004, 10'd201 }; 
        'd2196: dout <= { 2'd1, 8'd037, 10'd340 }; 
        'd2197: dout <= { 2'd1, 8'd015, 10'd074 }; 
        'd2198: dout <= { 2'd2, 8'd011, 10'd119 }; 
        'd2199: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd2200: dout <= { 2'd1, 8'd037, 10'd329 }; 
        'd2201: dout <= { 2'd1, 8'd003, 10'd103 }; 
        'd2202: dout <= { 2'd1, 8'd012, 10'd166 }; 
        'd2203: dout <= { 2'd1, 8'd016, 10'd242 }; 
        'd2204: dout <= { 2'd1, 8'd022, 10'd136 }; 
        'd2205: dout <= { 2'd1, 8'd049, 10'd295 }; 
        'd2206: dout <= { 2'd1, 8'd001, 10'd189 }; 
        'd2207: dout <= { 2'd1, 8'd036, 10'd092 }; 
        'd2208: dout <= { 2'd1, 8'd059, 10'd072 }; 
        'd2209: dout <= { 2'd1, 8'd034, 10'd290 }; 
        'd2210: dout <= { 2'd1, 8'd057, 10'd257 }; 
        'd2211: dout <= { 2'd2, 8'd052, 10'd308 }; 
        'd2212: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd2213: dout <= { 2'd1, 8'd031, 10'd077 }; 
        'd2214: dout <= { 2'd1, 8'd009, 10'd328 }; 
        'd2215: dout <= { 2'd1, 8'd048, 10'd026 }; 
        'd2216: dout <= { 2'd1, 8'd059, 10'd010 }; 
        'd2217: dout <= { 2'd1, 8'd027, 10'd278 }; 
        'd2218: dout <= { 2'd1, 8'd055, 10'd238 }; 
        'd2219: dout <= { 2'd1, 8'd023, 10'd102 }; 
        'd2220: dout <= { 2'd1, 8'd058, 10'd050 }; 
        'd2221: dout <= { 2'd1, 8'd038, 10'd243 }; 
        'd2222: dout <= { 2'd1, 8'd014, 10'd298 }; 
        'd2223: dout <= { 2'd1, 8'd044, 10'd344 }; 
        'd2224: dout <= { 2'd2, 8'd026, 10'd088 }; 
        'd2225: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd2226: dout <= { 2'd1, 8'd058, 10'd162 }; 
        'd2227: dout <= { 2'd1, 8'd032, 10'd042 }; 
        'd2228: dout <= { 2'd1, 8'd036, 10'd201 }; 
        'd2229: dout <= { 2'd1, 8'd009, 10'd206 }; 
        'd2230: dout <= { 2'd1, 8'd018, 10'd253 }; 
        'd2231: dout <= { 2'd1, 8'd030, 10'd281 }; 
        'd2232: dout <= { 2'd1, 8'd051, 10'd080 }; 
        'd2233: dout <= { 2'd1, 8'd049, 10'd051 }; 
        'd2234: dout <= { 2'd1, 8'd020, 10'd028 }; 
        'd2235: dout <= { 2'd1, 8'd005, 10'd312 }; 
        'd2236: dout <= { 2'd1, 8'd017, 10'd033 }; 
        'd2237: dout <= { 2'd2, 8'd042, 10'd264 }; 
        'd2238: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd2239: dout <= { 2'd1, 8'd006, 10'd008 }; 
        'd2240: dout <= { 2'd1, 8'd051, 10'd101 }; 
        'd2241: dout <= { 2'd1, 8'd003, 10'd229 }; 
        'd2242: dout <= { 2'd1, 8'd017, 10'd192 }; 
        'd2243: dout <= { 2'd1, 8'd011, 10'd093 }; 
        'd2244: dout <= { 2'd1, 8'd053, 10'd123 }; 
        'd2245: dout <= { 2'd1, 8'd047, 10'd253 }; 
        'd2246: dout <= { 2'd1, 8'd045, 10'd235 }; 
        'd2247: dout <= { 2'd1, 8'd043, 10'd024 }; 
        'd2248: dout <= { 2'd1, 8'd047, 10'd064 }; 
        'd2249: dout <= { 2'd1, 8'd031, 10'd290 }; 
        'd2250: dout <= { 2'd2, 8'd010, 10'd207 }; 
        'd2251: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd2252: dout <= { 2'd1, 8'd007, 10'd344 }; 
        'd2253: dout <= { 2'd1, 8'd031, 10'd238 }; 
        'd2254: dout <= { 2'd1, 8'd034, 10'd195 }; 
        'd2255: dout <= { 2'd1, 8'd040, 10'd069 }; 
        'd2256: dout <= { 2'd1, 8'd010, 10'd135 }; 
        'd2257: dout <= { 2'd1, 8'd005, 10'd092 }; 
        'd2258: dout <= { 2'd1, 8'd021, 10'd202 }; 
        'd2259: dout <= { 2'd1, 8'd041, 10'd262 }; 
        'd2260: dout <= { 2'd1, 8'd001, 10'd311 }; 
        'd2261: dout <= { 2'd1, 8'd021, 10'd307 }; 
        'd2262: dout <= { 2'd1, 8'd009, 10'd176 }; 
        'd2263: dout <= { 2'd2, 8'd032, 10'd136 }; 
        'd2264: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd2265: dout <= { 2'd1, 8'd011, 10'd063 }; 
        'd2266: dout <= { 2'd1, 8'd059, 10'd245 }; 
        'd2267: dout <= { 2'd1, 8'd024, 10'd254 }; 
        'd2268: dout <= { 2'd1, 8'd058, 10'd331 }; 
        'd2269: dout <= { 2'd1, 8'd052, 10'd168 }; 
        'd2270: dout <= { 2'd1, 8'd002, 10'd151 }; 
        'd2271: dout <= { 2'd1, 8'd050, 10'd166 }; 
        'd2272: dout <= { 2'd1, 8'd006, 10'd213 }; 
        'd2273: dout <= { 2'd1, 8'd055, 10'd177 }; 
        'd2274: dout <= { 2'd1, 8'd022, 10'd161 }; 
        'd2275: dout <= { 2'd1, 8'd046, 10'd320 }; 
        'd2276: dout <= { 2'd2, 8'd054, 10'd090 }; 
        'd2277: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd2278: dout <= { 2'd1, 8'd025, 10'd325 }; 
        'd2279: dout <= { 2'd1, 8'd005, 10'd158 }; 
        'd2280: dout <= { 2'd1, 8'd037, 10'd129 }; 
        'd2281: dout <= { 2'd1, 8'd019, 10'd333 }; 
        'd2282: dout <= { 2'd1, 8'd038, 10'd139 }; 
        'd2283: dout <= { 2'd1, 8'd029, 10'd153 }; 
        'd2284: dout <= { 2'd1, 8'd043, 10'd052 }; 
        'd2285: dout <= { 2'd1, 8'd012, 10'd337 }; 
        'd2286: dout <= { 2'd1, 8'd030, 10'd111 }; 
        'd2287: dout <= { 2'd1, 8'd018, 10'd275 }; 
        'd2288: dout <= { 2'd1, 8'd056, 10'd011 }; 
        'd2289: dout <= { 2'd2, 8'd033, 10'd122 }; 
        'd2290: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd2291: dout <= { 2'd1, 8'd028, 10'd076 }; 
        'd2292: dout <= { 2'd1, 8'd049, 10'd111 }; 
        'd2293: dout <= { 2'd1, 8'd042, 10'd336 }; 
        'd2294: dout <= { 2'd1, 8'd045, 10'd181 }; 
        'd2295: dout <= { 2'd1, 8'd015, 10'd015 }; 
        'd2296: dout <= { 2'd1, 8'd057, 10'd071 }; 
        'd2297: dout <= { 2'd1, 8'd033, 10'd184 }; 
        'd2298: dout <= { 2'd1, 8'd016, 10'd226 }; 
        'd2299: dout <= { 2'd1, 8'd053, 10'd273 }; 
        'd2300: dout <= { 2'd1, 8'd008, 10'd006 }; 
        'd2301: dout <= { 2'd1, 8'd028, 10'd058 }; 
        'd2302: dout <= { 2'd2, 8'd051, 10'd352 }; 
        'd2303: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd2304: dout <= { 2'd1, 8'd032, 10'd234 }; 
        'd2305: dout <= { 2'd1, 8'd013, 10'd067 }; 
        'd2306: dout <= { 2'd1, 8'd039, 10'd332 }; 
        'd2307: dout <= { 2'd1, 8'd008, 10'd210 }; 
        'd2308: dout <= { 2'd1, 8'd031, 10'd010 }; 
        'd2309: dout <= { 2'd1, 8'd054, 10'd324 }; 
        'd2310: dout <= { 2'd1, 8'd000, 10'd236 }; 
        'd2311: dout <= { 2'd1, 8'd029, 10'd137 }; 
        'd2312: dout <= { 2'd1, 8'd023, 10'd170 }; 
        'd2313: dout <= { 2'd1, 8'd024, 10'd358 }; 
        'd2314: dout <= { 2'd1, 8'd035, 10'd206 }; 
        'd2315: dout <= { 2'd2, 8'd002, 10'd072 }; 
        'd2316: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd2317: dout <= { 2'd1, 8'd000, 10'd230 }; 
        'd2318: dout <= { 2'd2, 8'd001, 10'd236 }; 
        'd2319: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd2320: dout <= { 2'd1, 8'd008, 10'd049 }; 
        'd2321: dout <= { 2'd2, 8'd047, 10'd160 }; 
        'd2322: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd2323: dout <= { 2'd1, 8'd053, 10'd244 }; 
        'd2324: dout <= { 2'd2, 8'd007, 10'd267 }; 
        'd2325: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd2326: dout <= { 2'd1, 8'd046, 10'd341 }; 
        'd2327: dout <= { 2'd2, 8'd042, 10'd184 }; 
        'd2328: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd2329: dout <= { 2'd1, 8'd003, 10'd019 }; 
        'd2330: dout <= { 2'd2, 8'd020, 10'd150 }; 
        'd2331: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd2332: dout <= { 2'd1, 8'd001, 10'd225 }; 
        'd2333: dout <= { 2'd2, 8'd054, 10'd066 }; 
        'd2334: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd2335: dout <= { 2'd1, 8'd048, 10'd025 }; 
        'd2336: dout <= { 2'd2, 8'd030, 10'd036 }; 
        'd2337: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd2338: dout <= { 2'd1, 8'd036, 10'd203 }; 
        'd2339: dout <= { 2'd2, 8'd016, 10'd359 }; 
        'd2340: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd2341: dout <= { 2'd1, 8'd055, 10'd034 }; 
        'd2342: dout <= { 2'd2, 8'd037, 10'd331 }; 
        'd2343: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd2344: dout <= { 2'd1, 8'd049, 10'd069 }; 
        'd2345: dout <= { 2'd2, 8'd038, 10'd132 }; 
        'd2346: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd2347: dout <= { 2'd1, 8'd040, 10'd265 }; 
        'd2348: dout <= { 2'd2, 8'd028, 10'd167 }; 
        'd2349: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd2350: dout <= { 2'd1, 8'd035, 10'd008 }; 
        'd2351: dout <= { 2'd2, 8'd014, 10'd210 }; 
        'd2352: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd2353: dout <= { 2'd1, 8'd041, 10'd141 }; 
        'd2354: dout <= { 2'd2, 8'd050, 10'd140 }; 
        'd2355: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd2356: dout <= { 2'd1, 8'd015, 10'd293 }; 
        'd2357: dout <= { 2'd2, 8'd044, 10'd279 }; 
        'd2358: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd2359: dout <= { 2'd1, 8'd033, 10'd098 }; 
        'd2360: dout <= { 2'd2, 8'd035, 10'd141 }; 
        'd2361: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd2362: dout <= { 2'd1, 8'd014, 10'd273 }; 
        'd2363: dout <= { 2'd2, 8'd043, 10'd173 }; 
        'd2364: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd2365: dout <= { 2'd1, 8'd029, 10'd123 }; 
        'd2366: dout <= { 2'd2, 8'd021, 10'd116 }; 
        'd2367: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd2368: dout <= { 2'd1, 8'd018, 10'd111 }; 
        'd2369: dout <= { 2'd2, 8'd039, 10'd265 }; 
        'd2370: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd2371: dout <= { 2'd1, 8'd004, 10'd339 }; 
        'd2372: dout <= { 2'd2, 8'd027, 10'd216 }; 
        'd2373: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd2374: dout <= { 2'd1, 8'd050, 10'd041 }; 
        'd2375: dout <= { 2'd2, 8'd008, 10'd243 }; 
        'd2376: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd2377: dout <= { 2'd1, 8'd038, 10'd298 }; 
        'd2378: dout <= { 2'd2, 8'd055, 10'd110 }; 
        'd2379: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd2380: dout <= { 2'd1, 8'd043, 10'd111 }; 
        'd2381: dout <= { 2'd2, 8'd011, 10'd324 }; 
        'd2382: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd2383: dout <= { 2'd1, 8'd016, 10'd008 }; 
        'd2384: dout <= { 2'd2, 8'd017, 10'd070 }; 
        'd2385: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd2386: dout <= { 2'd1, 8'd030, 10'd121 }; 
        'd2387: dout <= { 2'd2, 8'd006, 10'd096 }; 
        'd2388: dout <= { 2'd1, 8'd036, 10'd000 }; 
        'd2389: dout <= { 2'd1, 8'd021, 10'd175 }; 
        'd2390: dout <= { 2'd2, 8'd045, 10'd148 }; 
        'd2391: dout <= { 2'd1, 8'd037, 10'd000 }; 
        'd2392: dout <= { 2'd1, 8'd039, 10'd339 }; 
        'd2393: dout <= { 2'd2, 8'd025, 10'd198 }; 
        'd2394: dout <= { 2'd1, 8'd038, 10'd000 }; 
        'd2395: dout <= { 2'd1, 8'd010, 10'd068 }; 
        'd2396: dout <= { 2'd2, 8'd018, 10'd097 }; 
        'd2397: dout <= { 2'd1, 8'd039, 10'd000 }; 
        'd2398: dout <= { 2'd1, 8'd002, 10'd318 }; 
        'd2399: dout <= { 2'd2, 8'd000, 10'd284 }; 
        'd2400: dout <= { 2'd1, 8'd040, 10'd000 }; 
        'd2401: dout <= { 2'd1, 8'd013, 10'd337 }; 
        'd2402: dout <= { 2'd2, 8'd052, 10'd205 }; 
        'd2403: dout <= { 2'd1, 8'd041, 10'd000 }; 
        'd2404: dout <= { 2'd1, 8'd045, 10'd322 }; 
        'd2405: dout <= { 2'd2, 8'd046, 10'd325 }; 
        'd2406: dout <= { 2'd1, 8'd042, 10'd000 }; 
        'd2407: dout <= { 2'd1, 8'd009, 10'd104 }; 
        'd2408: dout <= { 2'd2, 8'd010, 10'd317 }; 
        'd2409: dout <= { 2'd1, 8'd043, 10'd000 }; 
        'd2410: dout <= { 2'd1, 8'd057, 10'd183 }; 
        'd2411: dout <= { 2'd2, 8'd053, 10'd319 }; 
        'd2412: dout <= { 2'd1, 8'd044, 10'd000 }; 
        'd2413: dout <= { 2'd1, 8'd020, 10'd329 }; 
        'd2414: dout <= { 2'd2, 8'd012, 10'd196 }; 
        'd2415: dout <= { 2'd1, 8'd045, 10'd000 }; 
        'd2416: dout <= { 2'd1, 8'd024, 10'd327 }; 
        'd2417: dout <= { 2'd2, 8'd048, 10'd123 }; 
        'd2418: dout <= { 2'd1, 8'd046, 10'd000 }; 
        'd2419: dout <= { 2'd1, 8'd056, 10'd267 }; 
        'd2420: dout <= { 2'd2, 8'd041, 10'd058 }; 
        'd2421: dout <= { 2'd1, 8'd047, 10'd000 }; 
        'd2422: dout <= { 2'd1, 8'd019, 10'd196 }; 
        'd2423: dout <= { 2'd2, 8'd002, 10'd351 }; 
        'd2424: dout <= { 2'd1, 8'd048, 10'd000 }; 
        'd2425: dout <= { 2'd1, 8'd042, 10'd217 }; 
        'd2426: dout <= { 2'd2, 8'd022, 10'd161 }; 
        'd2427: dout <= { 2'd1, 8'd049, 10'd000 }; 
        'd2428: dout <= { 2'd1, 8'd054, 10'd148 }; 
        'd2429: dout <= { 2'd2, 8'd057, 10'd086 }; 
        'd2430: dout <= { 2'd1, 8'd050, 10'd000 }; 
        'd2431: dout <= { 2'd1, 8'd047, 10'd184 }; 
        'd2432: dout <= { 2'd2, 8'd019, 10'd055 }; 
        'd2433: dout <= { 2'd1, 8'd051, 10'd000 }; 
        'd2434: dout <= { 2'd1, 8'd052, 10'd314 }; 
        'd2435: dout <= { 2'd2, 8'd036, 10'd072 }; 
        'd2436: dout <= { 2'd1, 8'd052, 10'd000 }; 
        'd2437: dout <= { 2'd1, 8'd034, 10'd131 }; 
        'd2438: dout <= { 2'd2, 8'd058, 10'd064 }; 
        'd2439: dout <= { 2'd1, 8'd053, 10'd000 }; 
        'd2440: dout <= { 2'd1, 8'd023, 10'd099 }; 
        'd2441: dout <= { 2'd2, 8'd040, 10'd072 }; 
        'd2442: dout <= { 2'd1, 8'd054, 10'd000 }; 
        'd2443: dout <= { 2'd1, 8'd026, 10'd122 }; 
        'd2444: dout <= { 2'd2, 8'd026, 10'd195 }; 
        'd2445: dout <= { 2'd1, 8'd055, 10'd000 }; 
        'd2446: dout <= { 2'd1, 8'd022, 10'd086 }; 
        'd2447: dout <= { 2'd2, 8'd029, 10'd093 }; 
        'd2448: dout <= { 2'd1, 8'd056, 10'd000 }; 
        'd2449: dout <= { 2'd1, 8'd012, 10'd040 }; 
        'd2450: dout <= { 2'd2, 8'd015, 10'd288 }; 
        'd2451: dout <= { 2'd1, 8'd057, 10'd000 }; 
        'd2452: dout <= { 2'd1, 8'd005, 10'd164 }; 
        'd2453: dout <= { 2'd2, 8'd034, 10'd341 }; 
        'd2454: dout <= { 2'd1, 8'd058, 10'd000 }; 
        'd2455: dout <= { 2'd1, 8'd027, 10'd111 }; 
        'd2456: dout <= { 2'd2, 8'd004, 10'd031 }; 
        'd2457: dout <= { 2'd1, 8'd059, 10'd000 }; 
        'd2458: dout <= { 2'd1, 8'd044, 10'd342 }; 
        'd2459: dout <= { 2'd2, 8'd056, 10'd086 }; 
        'd2460: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd2461: dout <= { 2'd1, 8'd046, 10'd303 }; 
        'd2462: dout <= { 2'd2, 8'd047, 10'd286 }; 
        'd2463: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd2464: dout <= { 2'd1, 8'd020, 10'd156 }; 
        'd2465: dout <= { 2'd2, 8'd046, 10'd137 }; 
        'd2466: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd2467: dout <= { 2'd1, 8'd053, 10'd117 }; 
        'd2468: dout <= { 2'd2, 8'd005, 10'd051 }; 
        'd2469: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd2470: dout <= { 2'd1, 8'd012, 10'd304 }; 
        'd2471: dout <= { 2'd2, 8'd057, 10'd223 }; 
        'd2472: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd2473: dout <= { 2'd1, 8'd041, 10'd152 }; 
        'd2474: dout <= { 2'd2, 8'd042, 10'd260 }; 
        'd2475: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd2476: dout <= { 2'd1, 8'd034, 10'd178 }; 
        'd2477: dout <= { 2'd2, 8'd013, 10'd169 }; 
        'd2478: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd2479: dout <= { 2'd1, 8'd005, 10'd193 }; 
        'd2480: dout <= { 2'd2, 8'd018, 10'd151 }; 
        'd2481: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd2482: dout <= { 2'd1, 8'd019, 10'd089 }; 
        'd2483: dout <= { 2'd2, 8'd058, 10'd156 }; 
        'd2484: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd2485: dout <= { 2'd1, 8'd024, 10'd150 }; 
        'd2486: dout <= { 2'd2, 8'd035, 10'd158 }; 
        'd2487: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd2488: dout <= { 2'd1, 8'd006, 10'd020 }; 
        'd2489: dout <= { 2'd2, 8'd034, 10'd272 }; 
        'd2490: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd2491: dout <= { 2'd1, 8'd054, 10'd249 }; 
        'd2492: dout <= { 2'd2, 8'd022, 10'd018 }; 
        'd2493: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd2494: dout <= { 2'd1, 8'd015, 10'd156 }; 
        'd2495: dout <= { 2'd2, 8'd036, 10'd346 }; 
        'd2496: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd2497: dout <= { 2'd1, 8'd004, 10'd266 }; 
        'd2498: dout <= { 2'd2, 8'd027, 10'd100 }; 
        'd2499: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd2500: dout <= { 2'd1, 8'd029, 10'd246 }; 
        'd2501: dout <= { 2'd2, 8'd032, 10'd107 }; 
        'd2502: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd2503: dout <= { 2'd1, 8'd022, 10'd133 }; 
        'd2504: dout <= { 2'd2, 8'd051, 10'd309 }; 
        'd2505: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd2506: dout <= { 2'd1, 8'd042, 10'd245 }; 
        'd2507: dout <= { 2'd2, 8'd049, 10'd234 }; 
        'd2508: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd2509: dout <= { 2'd1, 8'd013, 10'd004 }; 
        'd2510: dout <= { 2'd2, 8'd045, 10'd050 }; 
        'd2511: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd2512: dout <= { 2'd1, 8'd014, 10'd021 }; 
        'd2513: dout <= { 2'd2, 8'd026, 10'd321 }; 
        'd2514: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd2515: dout <= { 2'd1, 8'd017, 10'd246 }; 
        'd2516: dout <= { 2'd2, 8'd004, 10'd034 }; 
        'd2517: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd2518: dout <= { 2'd1, 8'd000, 10'd232 }; 
        'd2519: dout <= { 2'd2, 8'd000, 10'd165 }; 
        'd2520: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd2521: dout <= { 2'd1, 8'd032, 10'd007 }; 
        'd2522: dout <= { 2'd2, 8'd054, 10'd122 }; 
        'd2523: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd2524: dout <= { 2'd1, 8'd026, 10'd303 }; 
        'd2525: dout <= { 2'd2, 8'd021, 10'd165 }; 
        'd2526: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd2527: dout <= { 2'd1, 8'd011, 10'd102 }; 
        'd2528: dout <= { 2'd2, 8'd014, 10'd090 }; 
        'd2529: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd2530: dout <= { 2'd1, 8'd057, 10'd167 }; 
        'd2531: dout <= { 2'd2, 8'd006, 10'd162 }; 
        'd2532: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd2533: dout <= { 2'd1, 8'd045, 10'd200 }; 
        'd2534: dout <= { 2'd2, 8'd019, 10'd091 }; 
        'd2535: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd2536: dout <= { 2'd1, 8'd002, 10'd072 }; 
        'd2537: dout <= { 2'd2, 8'd010, 10'd133 }; 
        'd2538: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd2539: dout <= { 2'd1, 8'd016, 10'd260 }; 
        'd2540: dout <= { 2'd2, 8'd030, 10'd092 }; 
        'd2541: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd2542: dout <= { 2'd1, 8'd021, 10'd259 }; 
        'd2543: dout <= { 2'd2, 8'd041, 10'd177 }; 
        'd2544: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd2545: dout <= { 2'd1, 8'd018, 10'd345 }; 
        'd2546: dout <= { 2'd2, 8'd007, 10'd123 }; 
        'd2547: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd2548: dout <= { 2'd1, 8'd058, 10'd041 }; 
        'd2549: dout <= { 2'd2, 8'd024, 10'd313 }; 
        'd2550: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd2551: dout <= { 2'd1, 8'd044, 10'd149 }; 
        'd2552: dout <= { 2'd2, 8'd020, 10'd043 }; 
        'd2553: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd2554: dout <= { 2'd1, 8'd036, 10'd108 }; 
        'd2555: dout <= { 2'd2, 8'd029, 10'd298 }; 
        'd2556: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd2557: dout <= { 2'd1, 8'd048, 10'd185 }; 
        'd2558: dout <= { 2'd2, 8'd038, 10'd001 }; 
        'd2559: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd2560: dout <= { 2'd1, 8'd039, 10'd342 }; 
        'd2561: dout <= { 2'd2, 8'd044, 10'd061 }; 
        'd2562: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd2563: dout <= { 2'd1, 8'd010, 10'd125 }; 
        'd2564: dout <= { 2'd2, 8'd009, 10'd026 }; 
        'd2565: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd2566: dout <= { 2'd1, 8'd040, 10'd266 }; 
        'd2567: dout <= { 2'd2, 8'd052, 10'd194 }; 
        'd2568: dout <= { 2'd1, 8'd036, 10'd000 }; 
        'd2569: dout <= { 2'd1, 8'd027, 10'd152 }; 
        'd2570: dout <= { 2'd2, 8'd043, 10'd171 }; 
        'd2571: dout <= { 2'd1, 8'd037, 10'd000 }; 
        'd2572: dout <= { 2'd1, 8'd030, 10'd277 }; 
        'd2573: dout <= { 2'd2, 8'd011, 10'd003 }; 
        'd2574: dout <= { 2'd1, 8'd038, 10'd000 }; 
        'd2575: dout <= { 2'd1, 8'd037, 10'd259 }; 
        'd2576: dout <= { 2'd2, 8'd025, 10'd311 }; 
        'd2577: dout <= { 2'd1, 8'd039, 10'd000 }; 
        'd2578: dout <= { 2'd1, 8'd007, 10'd286 }; 
        'd2579: dout <= { 2'd2, 8'd037, 10'd348 }; 
        'd2580: dout <= { 2'd1, 8'd040, 10'd000 }; 
        'd2581: dout <= { 2'd1, 8'd056, 10'd070 }; 
        'd2582: dout <= { 2'd2, 8'd031, 10'd056 }; 
        'd2583: dout <= { 2'd1, 8'd041, 10'd000 }; 
        'd2584: dout <= { 2'd1, 8'd052, 10'd334 }; 
        'd2585: dout <= { 2'd2, 8'd059, 10'd286 }; 
        'd2586: dout <= { 2'd1, 8'd042, 10'd000 }; 
        'd2587: dout <= { 2'd1, 8'd038, 10'd153 }; 
        'd2588: dout <= { 2'd2, 8'd016, 10'd084 }; 
        'd2589: dout <= { 2'd1, 8'd043, 10'd000 }; 
        'd2590: dout <= { 2'd1, 8'd009, 10'd307 }; 
        'd2591: dout <= { 2'd2, 8'd012, 10'd141 }; 
        'd2592: dout <= { 2'd1, 8'd044, 10'd000 }; 
        'd2593: dout <= { 2'd1, 8'd033, 10'd201 }; 
        'd2594: dout <= { 2'd2, 8'd053, 10'd345 }; 
        'd2595: dout <= { 2'd1, 8'd045, 10'd000 }; 
        'd2596: dout <= { 2'd1, 8'd025, 10'd272 }; 
        'd2597: dout <= { 2'd2, 8'd028, 10'd212 }; 
        'd2598: dout <= { 2'd1, 8'd046, 10'd000 }; 
        'd2599: dout <= { 2'd1, 8'd003, 10'd267 }; 
        'd2600: dout <= { 2'd2, 8'd055, 10'd184 }; 
        'd2601: dout <= { 2'd1, 8'd047, 10'd000 }; 
        'd2602: dout <= { 2'd1, 8'd008, 10'd084 }; 
        'd2603: dout <= { 2'd2, 8'd015, 10'd293 }; 
        'd2604: dout <= { 2'd1, 8'd048, 10'd000 }; 
        'd2605: dout <= { 2'd1, 8'd035, 10'd316 }; 
        'd2606: dout <= { 2'd2, 8'd017, 10'd080 }; 
        'd2607: dout <= { 2'd1, 8'd049, 10'd000 }; 
        'd2608: dout <= { 2'd1, 8'd043, 10'd274 }; 
        'd2609: dout <= { 2'd2, 8'd056, 10'd058 }; 
        'd2610: dout <= { 2'd1, 8'd050, 10'd000 }; 
        'd2611: dout <= { 2'd1, 8'd059, 10'd023 }; 
        'd2612: dout <= { 2'd2, 8'd008, 10'd269 }; 
        'd2613: dout <= { 2'd1, 8'd051, 10'd000 }; 
        'd2614: dout <= { 2'd1, 8'd001, 10'd061 }; 
        'd2615: dout <= { 2'd2, 8'd039, 10'd050 }; 
        'd2616: dout <= { 2'd1, 8'd052, 10'd000 }; 
        'd2617: dout <= { 2'd1, 8'd050, 10'd316 }; 
        'd2618: dout <= { 2'd2, 8'd001, 10'd302 }; 
        'd2619: dout <= { 2'd1, 8'd053, 10'd000 }; 
        'd2620: dout <= { 2'd1, 8'd028, 10'd149 }; 
        'd2621: dout <= { 2'd2, 8'd033, 10'd196 }; 
        'd2622: dout <= { 2'd1, 8'd054, 10'd000 }; 
        'd2623: dout <= { 2'd1, 8'd047, 10'd223 }; 
        'd2624: dout <= { 2'd2, 8'd003, 10'd300 }; 
        'd2625: dout <= { 2'd1, 8'd055, 10'd000 }; 
        'd2626: dout <= { 2'd1, 8'd023, 10'd088 }; 
        'd2627: dout <= { 2'd2, 8'd023, 10'd051 }; 
        'd2628: dout <= { 2'd1, 8'd056, 10'd000 }; 
        'd2629: dout <= { 2'd1, 8'd051, 10'd008 }; 
        'd2630: dout <= { 2'd2, 8'd048, 10'd277 }; 
        'd2631: dout <= { 2'd1, 8'd057, 10'd000 }; 
        'd2632: dout <= { 2'd1, 8'd031, 10'd079 }; 
        'd2633: dout <= { 2'd2, 8'd002, 10'd112 }; 
        'd2634: dout <= { 2'd1, 8'd058, 10'd000 }; 
        'd2635: dout <= { 2'd1, 8'd055, 10'd094 }; 
        'd2636: dout <= { 2'd2, 8'd040, 10'd132 }; 
        'd2637: dout <= { 2'd1, 8'd059, 10'd000 }; 
        'd2638: dout <= { 2'd1, 8'd049, 10'd059 }; 
        'd2639: dout <= { 2'd3, 8'd050, 10'd243 }; 
        // Q=45, BaseAddr=2640
        'd2640: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd2641: dout <= { 2'd1, 8'd040, 10'd141 }; 
        'd2642: dout <= { 2'd1, 8'd026, 10'd175 }; 
        'd2643: dout <= { 2'd1, 8'd031, 10'd324 }; 
        'd2644: dout <= { 2'd1, 8'd024, 10'd297 }; 
        'd2645: dout <= { 2'd1, 8'd040, 10'd248 }; 
        'd2646: dout <= { 2'd1, 8'd012, 10'd072 }; 
        'd2647: dout <= { 2'd1, 8'd023, 10'd116 }; 
        'd2648: dout <= { 2'd1, 8'd029, 10'd055 }; 
        'd2649: dout <= { 2'd1, 8'd022, 10'd060 }; 
        'd2650: dout <= { 2'd1, 8'd011, 10'd018 }; 
        'd2651: dout <= { 2'd2, 8'd039, 10'd163 }; 
        'd2652: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd2653: dout <= { 2'd1, 8'd019, 10'd252 }; 
        'd2654: dout <= { 2'd1, 8'd043, 10'd059 }; 
        'd2655: dout <= { 2'd1, 8'd042, 10'd007 }; 
        'd2656: dout <= { 2'd1, 8'd009, 10'd307 }; 
        'd2657: dout <= { 2'd1, 8'd037, 10'd283 }; 
        'd2658: dout <= { 2'd1, 8'd044, 10'd160 }; 
        'd2659: dout <= { 2'd1, 8'd002, 10'd150 }; 
        'd2660: dout <= { 2'd1, 8'd010, 10'd340 }; 
        'd2661: dout <= { 2'd1, 8'd042, 10'd018 }; 
        'd2662: dout <= { 2'd1, 8'd021, 10'd044 }; 
        'd2663: dout <= { 2'd2, 8'd032, 10'd253 }; 
        'd2664: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd2665: dout <= { 2'd1, 8'd032, 10'd174 }; 
        'd2666: dout <= { 2'd1, 8'd012, 10'd177 }; 
        'd2667: dout <= { 2'd1, 8'd021, 10'd140 }; 
        'd2668: dout <= { 2'd1, 8'd022, 10'd302 }; 
        'd2669: dout <= { 2'd1, 8'd002, 10'd271 }; 
        'd2670: dout <= { 2'd1, 8'd004, 10'd321 }; 
        'd2671: dout <= { 2'd1, 8'd017, 10'd336 }; 
        'd2672: dout <= { 2'd1, 8'd000, 10'd308 }; 
        'd2673: dout <= { 2'd1, 8'd043, 10'd037 }; 
        'd2674: dout <= { 2'd1, 8'd009, 10'd142 }; 
        'd2675: dout <= { 2'd2, 8'd034, 10'd298 }; 
        'd2676: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd2677: dout <= { 2'd1, 8'd030, 10'd034 }; 
        'd2678: dout <= { 2'd1, 8'd014, 10'd262 }; 
        'd2679: dout <= { 2'd1, 8'd000, 10'd155 }; 
        'd2680: dout <= { 2'd1, 8'd017, 10'd295 }; 
        'd2681: dout <= { 2'd1, 8'd001, 10'd081 }; 
        'd2682: dout <= { 2'd1, 8'd032, 10'd084 }; 
        'd2683: dout <= { 2'd1, 8'd042, 10'd194 }; 
        'd2684: dout <= { 2'd1, 8'd016, 10'd162 }; 
        'd2685: dout <= { 2'd1, 8'd035, 10'd128 }; 
        'd2686: dout <= { 2'd1, 8'd017, 10'd318 }; 
        'd2687: dout <= { 2'd2, 8'd036, 10'd174 }; 
        'd2688: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd2689: dout <= { 2'd1, 8'd021, 10'd169 }; 
        'd2690: dout <= { 2'd1, 8'd022, 10'd253 }; 
        'd2691: dout <= { 2'd1, 8'd019, 10'd324 }; 
        'd2692: dout <= { 2'd1, 8'd014, 10'd215 }; 
        'd2693: dout <= { 2'd1, 8'd008, 10'd036 }; 
        'd2694: dout <= { 2'd1, 8'd043, 10'd046 }; 
        'd2695: dout <= { 2'd1, 8'd009, 10'd240 }; 
        'd2696: dout <= { 2'd1, 8'd013, 10'd206 }; 
        'd2697: dout <= { 2'd1, 8'd015, 10'd027 }; 
        'd2698: dout <= { 2'd1, 8'd031, 10'd338 }; 
        'd2699: dout <= { 2'd2, 8'd010, 10'd108 }; 
        'd2700: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd2701: dout <= { 2'd1, 8'd035, 10'd035 }; 
        'd2702: dout <= { 2'd1, 8'd029, 10'd126 }; 
        'd2703: dout <= { 2'd1, 8'd036, 10'd352 }; 
        'd2704: dout <= { 2'd1, 8'd041, 10'd209 }; 
        'd2705: dout <= { 2'd1, 8'd005, 10'd278 }; 
        'd2706: dout <= { 2'd1, 8'd005, 10'd031 }; 
        'd2707: dout <= { 2'd1, 8'd003, 10'd140 }; 
        'd2708: dout <= { 2'd1, 8'd011, 10'd120 }; 
        'd2709: dout <= { 2'd1, 8'd006, 10'd315 }; 
        'd2710: dout <= { 2'd1, 8'd020, 10'd309 }; 
        'd2711: dout <= { 2'd2, 8'd023, 10'd163 }; 
        'd2712: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd2713: dout <= { 2'd1, 8'd009, 10'd090 }; 
        'd2714: dout <= { 2'd1, 8'd016, 10'd196 }; 
        'd2715: dout <= { 2'd1, 8'd030, 10'd075 }; 
        'd2716: dout <= { 2'd1, 8'd023, 10'd174 }; 
        'd2717: dout <= { 2'd1, 8'd027, 10'd177 }; 
        'd2718: dout <= { 2'd1, 8'd036, 10'd340 }; 
        'd2719: dout <= { 2'd1, 8'd030, 10'd132 }; 
        'd2720: dout <= { 2'd1, 8'd018, 10'd230 }; 
        'd2721: dout <= { 2'd1, 8'd018, 10'd228 }; 
        'd2722: dout <= { 2'd1, 8'd000, 10'd215 }; 
        'd2723: dout <= { 2'd2, 8'd016, 10'd103 }; 
        'd2724: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd2725: dout <= { 2'd1, 8'd031, 10'd098 }; 
        'd2726: dout <= { 2'd1, 8'd003, 10'd088 }; 
        'd2727: dout <= { 2'd1, 8'd018, 10'd203 }; 
        'd2728: dout <= { 2'd1, 8'd039, 10'd046 }; 
        'd2729: dout <= { 2'd1, 8'd038, 10'd281 }; 
        'd2730: dout <= { 2'd1, 8'd034, 10'd165 }; 
        'd2731: dout <= { 2'd1, 8'd015, 10'd267 }; 
        'd2732: dout <= { 2'd1, 8'd026, 10'd271 }; 
        'd2733: dout <= { 2'd1, 8'd044, 10'd013 }; 
        'd2734: dout <= { 2'd1, 8'd002, 10'd338 }; 
        'd2735: dout <= { 2'd2, 8'd001, 10'd009 }; 
        'd2736: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd2737: dout <= { 2'd1, 8'd022, 10'd133 }; 
        'd2738: dout <= { 2'd1, 8'd041, 10'd186 }; 
        'd2739: dout <= { 2'd1, 8'd011, 10'd128 }; 
        'd2740: dout <= { 2'd1, 8'd032, 10'd077 }; 
        'd2741: dout <= { 2'd1, 8'd003, 10'd012 }; 
        'd2742: dout <= { 2'd1, 8'd027, 10'd315 }; 
        'd2743: dout <= { 2'd1, 8'd020, 10'd019 }; 
        'd2744: dout <= { 2'd1, 8'd006, 10'd204 }; 
        'd2745: dout <= { 2'd1, 8'd025, 10'd138 }; 
        'd2746: dout <= { 2'd1, 8'd003, 10'd309 }; 
        'd2747: dout <= { 2'd2, 8'd008, 10'd079 }; 
        'd2748: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd2749: dout <= { 2'd1, 8'd037, 10'd071 }; 
        'd2750: dout <= { 2'd1, 8'd010, 10'd147 }; 
        'd2751: dout <= { 2'd1, 8'd025, 10'd106 }; 
        'd2752: dout <= { 2'd1, 8'd006, 10'd012 }; 
        'd2753: dout <= { 2'd1, 8'd016, 10'd217 }; 
        'd2754: dout <= { 2'd1, 8'd001, 10'd046 }; 
        'd2755: dout <= { 2'd1, 8'd022, 10'd162 }; 
        'd2756: dout <= { 2'd1, 8'd024, 10'd075 }; 
        'd2757: dout <= { 2'd1, 8'd005, 10'd161 }; 
        'd2758: dout <= { 2'd1, 8'd027, 10'd109 }; 
        'd2759: dout <= { 2'd2, 8'd007, 10'd281 }; 
        'd2760: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd2761: dout <= { 2'd1, 8'd000, 10'd196 }; 
        'd2762: dout <= { 2'd1, 8'd008, 10'd224 }; 
        'd2763: dout <= { 2'd1, 8'd020, 10'd246 }; 
        'd2764: dout <= { 2'd1, 8'd004, 10'd157 }; 
        'd2765: dout <= { 2'd1, 8'd015, 10'd146 }; 
        'd2766: dout <= { 2'd1, 8'd039, 10'd291 }; 
        'd2767: dout <= { 2'd1, 8'd033, 10'd225 }; 
        'd2768: dout <= { 2'd1, 8'd028, 10'd159 }; 
        'd2769: dout <= { 2'd1, 8'd038, 10'd010 }; 
        'd2770: dout <= { 2'd1, 8'd030, 10'd165 }; 
        'd2771: dout <= { 2'd2, 8'd013, 10'd205 }; 
        'd2772: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd2773: dout <= { 2'd1, 8'd013, 10'd042 }; 
        'd2774: dout <= { 2'd1, 8'd018, 10'd240 }; 
        'd2775: dout <= { 2'd1, 8'd029, 10'd002 }; 
        'd2776: dout <= { 2'd1, 8'd035, 10'd004 }; 
        'd2777: dout <= { 2'd1, 8'd043, 10'd167 }; 
        'd2778: dout <= { 2'd1, 8'd021, 10'd245 }; 
        'd2779: dout <= { 2'd1, 8'd040, 10'd235 }; 
        'd2780: dout <= { 2'd1, 8'd025, 10'd256 }; 
        'd2781: dout <= { 2'd1, 8'd024, 10'd328 }; 
        'd2782: dout <= { 2'd1, 8'd041, 10'd176 }; 
        'd2783: dout <= { 2'd2, 8'd004, 10'd347 }; 
        'd2784: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd2785: dout <= { 2'd1, 8'd010, 10'd081 }; 
        'd2786: dout <= { 2'd1, 8'd006, 10'd194 }; 
        'd2787: dout <= { 2'd1, 8'd012, 10'd109 }; 
        'd2788: dout <= { 2'd1, 8'd034, 10'd352 }; 
        'd2789: dout <= { 2'd1, 8'd044, 10'd113 }; 
        'd2790: dout <= { 2'd1, 8'd019, 10'd047 }; 
        'd2791: dout <= { 2'd1, 8'd014, 10'd354 }; 
        'd2792: dout <= { 2'd1, 8'd008, 10'd328 }; 
        'd2793: dout <= { 2'd1, 8'd040, 10'd158 }; 
        'd2794: dout <= { 2'd1, 8'd037, 10'd059 }; 
        'd2795: dout <= { 2'd2, 8'd029, 10'd032 }; 
        'd2796: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd2797: dout <= { 2'd1, 8'd036, 10'd184 }; 
        'd2798: dout <= { 2'd1, 8'd040, 10'd084 }; 
        'd2799: dout <= { 2'd1, 8'd010, 10'd011 }; 
        'd2800: dout <= { 2'd1, 8'd013, 10'd198 }; 
        'd2801: dout <= { 2'd1, 8'd007, 10'd150 }; 
        'd2802: dout <= { 2'd1, 8'd041, 10'd017 }; 
        'd2803: dout <= { 2'd1, 8'd037, 10'd176 }; 
        'd2804: dout <= { 2'd1, 8'd031, 10'd093 }; 
        'd2805: dout <= { 2'd1, 8'd019, 10'd346 }; 
        'd2806: dout <= { 2'd1, 8'd014, 10'd294 }; 
        'd2807: dout <= { 2'd2, 8'd012, 10'd058 }; 
        'd2808: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd2809: dout <= { 2'd1, 8'd018, 10'd321 }; 
        'd2810: dout <= { 2'd1, 8'd037, 10'd107 }; 
        'd2811: dout <= { 2'd1, 8'd028, 10'd349 }; 
        'd2812: dout <= { 2'd1, 8'd026, 10'd067 }; 
        'd2813: dout <= { 2'd1, 8'd033, 10'd248 }; 
        'd2814: dout <= { 2'd1, 8'd035, 10'd285 }; 
        'd2815: dout <= { 2'd1, 8'd038, 10'd303 }; 
        'd2816: dout <= { 2'd1, 8'd007, 10'd181 }; 
        'd2817: dout <= { 2'd1, 8'd026, 10'd145 }; 
        'd2818: dout <= { 2'd1, 8'd033, 10'd335 }; 
        'd2819: dout <= { 2'd2, 8'd028, 10'd194 }; 
        'd2820: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd2821: dout <= { 2'd1, 8'd044, 10'd069 }; 
        'd2822: dout <= { 2'd2, 8'd011, 10'd266 }; 
        'd2823: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd2824: dout <= { 2'd1, 8'd006, 10'd298 }; 
        'd2825: dout <= { 2'd2, 8'd021, 10'd153 }; 
        'd2826: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd2827: dout <= { 2'd1, 8'd003, 10'd291 }; 
        'd2828: dout <= { 2'd2, 8'd032, 10'd296 }; 
        'd2829: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd2830: dout <= { 2'd1, 8'd029, 10'd044 }; 
        'd2831: dout <= { 2'd2, 8'd015, 10'd321 }; 
        'd2832: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd2833: dout <= { 2'd1, 8'd007, 10'd160 }; 
        'd2834: dout <= { 2'd2, 8'd039, 10'd095 }; 
        'd2835: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd2836: dout <= { 2'd1, 8'd027, 10'd073 }; 
        'd2837: dout <= { 2'd2, 8'd030, 10'd087 }; 
        'd2838: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd2839: dout <= { 2'd1, 8'd008, 10'd098 }; 
        'd2840: dout <= { 2'd2, 8'd038, 10'd138 }; 
        'd2841: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd2842: dout <= { 2'd1, 8'd014, 10'd059 }; 
        'd2843: dout <= { 2'd2, 8'd025, 10'd310 }; 
        'd2844: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd2845: dout <= { 2'd1, 8'd011, 10'd168 }; 
        'd2846: dout <= { 2'd2, 8'd023, 10'd200 }; 
        'd2847: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd2848: dout <= { 2'd1, 8'd042, 10'd314 }; 
        'd2849: dout <= { 2'd2, 8'd042, 10'd065 }; 
        'd2850: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd2851: dout <= { 2'd1, 8'd026, 10'd161 }; 
        'd2852: dout <= { 2'd2, 8'd028, 10'd158 }; 
        'd2853: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd2854: dout <= { 2'd1, 8'd015, 10'd136 }; 
        'd2855: dout <= { 2'd2, 8'd035, 10'd303 }; 
        'd2856: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd2857: dout <= { 2'd1, 8'd020, 10'd166 }; 
        'd2858: dout <= { 2'd2, 8'd024, 10'd323 }; 
        'd2859: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd2860: dout <= { 2'd1, 8'd017, 10'd192 }; 
        'd2861: dout <= { 2'd2, 8'd036, 10'd054 }; 
        'd2862: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd2863: dout <= { 2'd1, 8'd004, 10'd191 }; 
        'd2864: dout <= { 2'd2, 8'd009, 10'd285 }; 
        'd2865: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd2866: dout <= { 2'd1, 8'd005, 10'd077 }; 
        'd2867: dout <= { 2'd2, 8'd002, 10'd070 }; 
        'd2868: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd2869: dout <= { 2'd1, 8'd012, 10'd309 }; 
        'd2870: dout <= { 2'd2, 8'd000, 10'd097 }; 
        'd2871: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd2872: dout <= { 2'd1, 8'd039, 10'd133 }; 
        'd2873: dout <= { 2'd2, 8'd005, 10'd305 }; 
        'd2874: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd2875: dout <= { 2'd1, 8'd038, 10'd243 }; 
        'd2876: dout <= { 2'd2, 8'd007, 10'd315 }; 
        'd2877: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd2878: dout <= { 2'd1, 8'd034, 10'd054 }; 
        'd2879: dout <= { 2'd2, 8'd027, 10'd292 }; 
        'd2880: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd2881: dout <= { 2'd1, 8'd016, 10'd117 }; 
        'd2882: dout <= { 2'd2, 8'd019, 10'd334 }; 
        'd2883: dout <= { 2'd1, 8'd036, 10'd000 }; 
        'd2884: dout <= { 2'd1, 8'd023, 10'd024 }; 
        'd2885: dout <= { 2'd2, 8'd004, 10'd041 }; 
        'd2886: dout <= { 2'd1, 8'd037, 10'd000 }; 
        'd2887: dout <= { 2'd1, 8'd033, 10'd045 }; 
        'd2888: dout <= { 2'd2, 8'd034, 10'd023 }; 
        'd2889: dout <= { 2'd1, 8'd038, 10'd000 }; 
        'd2890: dout <= { 2'd1, 8'd024, 10'd214 }; 
        'd2891: dout <= { 2'd2, 8'd020, 10'd135 }; 
        'd2892: dout <= { 2'd1, 8'd039, 10'd000 }; 
        'd2893: dout <= { 2'd1, 8'd001, 10'd318 }; 
        'd2894: dout <= { 2'd2, 8'd017, 10'd170 }; 
        'd2895: dout <= { 2'd1, 8'd040, 10'd000 }; 
        'd2896: dout <= { 2'd1, 8'd002, 10'd347 }; 
        'd2897: dout <= { 2'd2, 8'd001, 10'd181 }; 
        'd2898: dout <= { 2'd1, 8'd041, 10'd000 }; 
        'd2899: dout <= { 2'd1, 8'd043, 10'd101 }; 
        'd2900: dout <= { 2'd2, 8'd013, 10'd249 }; 
        'd2901: dout <= { 2'd1, 8'd042, 10'd000 }; 
        'd2902: dout <= { 2'd1, 8'd025, 10'd303 }; 
        'd2903: dout <= { 2'd2, 8'd033, 10'd138 }; 
        'd2904: dout <= { 2'd1, 8'd043, 10'd000 }; 
        'd2905: dout <= { 2'd1, 8'd028, 10'd190 }; 
        'd2906: dout <= { 2'd2, 8'd044, 10'd174 }; 
        'd2907: dout <= { 2'd1, 8'd044, 10'd000 }; 
        'd2908: dout <= { 2'd1, 8'd041, 10'd260 }; 
        'd2909: dout <= { 2'd2, 8'd031, 10'd059 }; 
        'd2910: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd2911: dout <= { 2'd1, 8'd032, 10'd022 }; 
        'd2912: dout <= { 2'd2, 8'd004, 10'd028 }; 
        'd2913: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd2914: dout <= { 2'd1, 8'd004, 10'd280 }; 
        'd2915: dout <= { 2'd2, 8'd020, 10'd221 }; 
        'd2916: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd2917: dout <= { 2'd1, 8'd027, 10'd182 }; 
        'd2918: dout <= { 2'd2, 8'd007, 10'd060 }; 
        'd2919: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd2920: dout <= { 2'd1, 8'd006, 10'd070 }; 
        'd2921: dout <= { 2'd2, 8'd003, 10'd262 }; 
        'd2922: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd2923: dout <= { 2'd1, 8'd039, 10'd007 }; 
        'd2924: dout <= { 2'd2, 8'd029, 10'd033 }; 
        'd2925: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd2926: dout <= { 2'd1, 8'd003, 10'd155 }; 
        'd2927: dout <= { 2'd2, 8'd018, 10'd312 }; 
        'd2928: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd2929: dout <= { 2'd1, 8'd002, 10'd176 }; 
        'd2930: dout <= { 2'd2, 8'd014, 10'd357 }; 
        'd2931: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd2932: dout <= { 2'd1, 8'd012, 10'd335 }; 
        'd2933: dout <= { 2'd2, 8'd033, 10'd269 }; 
        'd2934: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd2935: dout <= { 2'd1, 8'd013, 10'd112 }; 
        'd2936: dout <= { 2'd2, 8'd035, 10'd143 }; 
        'd2937: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd2938: dout <= { 2'd1, 8'd042, 10'd281 }; 
        'd2939: dout <= { 2'd2, 8'd037, 10'd331 }; 
        'd2940: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd2941: dout <= { 2'd1, 8'd023, 10'd343 }; 
        'd2942: dout <= { 2'd2, 8'd008, 10'd039 }; 
        'd2943: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd2944: dout <= { 2'd1, 8'd021, 10'd180 }; 
        'd2945: dout <= { 2'd2, 8'd011, 10'd038 }; 
        'd2946: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd2947: dout <= { 2'd1, 8'd011, 10'd276 }; 
        'd2948: dout <= { 2'd2, 8'd009, 10'd012 }; 
        'd2949: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd2950: dout <= { 2'd1, 8'd034, 10'd091 }; 
        'd2951: dout <= { 2'd2, 8'd026, 10'd157 }; 
        'd2952: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd2953: dout <= { 2'd1, 8'd031, 10'd031 }; 
        'd2954: dout <= { 2'd2, 8'd000, 10'd187 }; 
        'd2955: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd2956: dout <= { 2'd1, 8'd018, 10'd217 }; 
        'd2957: dout <= { 2'd2, 8'd044, 10'd168 }; 
        'd2958: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd2959: dout <= { 2'd1, 8'd040, 10'd139 }; 
        'd2960: dout <= { 2'd2, 8'd034, 10'd251 }; 
        'd2961: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd2962: dout <= { 2'd1, 8'd014, 10'd031 }; 
        'd2963: dout <= { 2'd2, 8'd001, 10'd268 }; 
        'd2964: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd2965: dout <= { 2'd1, 8'd010, 10'd179 }; 
        'd2966: dout <= { 2'd2, 8'd042, 10'd201 }; 
        'd2967: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd2968: dout <= { 2'd1, 8'd038, 10'd064 }; 
        'd2969: dout <= { 2'd2, 8'd023, 10'd187 }; 
        'd2970: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd2971: dout <= { 2'd1, 8'd033, 10'd028 }; 
        'd2972: dout <= { 2'd2, 8'd030, 10'd313 }; 
        'd2973: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd2974: dout <= { 2'd1, 8'd007, 10'd087 }; 
        'd2975: dout <= { 2'd2, 8'd036, 10'd307 }; 
        'd2976: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd2977: dout <= { 2'd1, 8'd026, 10'd085 }; 
        'd2978: dout <= { 2'd2, 8'd040, 10'd088 }; 
        'd2979: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd2980: dout <= { 2'd1, 8'd015, 10'd130 }; 
        'd2981: dout <= { 2'd2, 8'd013, 10'd039 }; 
        'd2982: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd2983: dout <= { 2'd1, 8'd000, 10'd059 }; 
        'd2984: dout <= { 2'd2, 8'd017, 10'd332 }; 
        'd2985: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd2986: dout <= { 2'd1, 8'd030, 10'd123 }; 
        'd2987: dout <= { 2'd2, 8'd032, 10'd140 }; 
        'd2988: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd2989: dout <= { 2'd1, 8'd028, 10'd095 }; 
        'd2990: dout <= { 2'd2, 8'd031, 10'd280 }; 
        'd2991: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd2992: dout <= { 2'd1, 8'd043, 10'd258 }; 
        'd2993: dout <= { 2'd2, 8'd041, 10'd271 }; 
        'd2994: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd2995: dout <= { 2'd1, 8'd005, 10'd356 }; 
        'd2996: dout <= { 2'd2, 8'd027, 10'd169 }; 
        'd2997: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd2998: dout <= { 2'd1, 8'd020, 10'd103 }; 
        'd2999: dout <= { 2'd2, 8'd043, 10'd313 }; 
        'd3000: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd3001: dout <= { 2'd1, 8'd044, 10'd212 }; 
        'd3002: dout <= { 2'd2, 8'd028, 10'd291 }; 
        'd3003: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd3004: dout <= { 2'd1, 8'd037, 10'd310 }; 
        'd3005: dout <= { 2'd2, 8'd012, 10'd213 }; 
        'd3006: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd3007: dout <= { 2'd1, 8'd019, 10'd342 }; 
        'd3008: dout <= { 2'd2, 8'd005, 10'd269 }; 
        'd3009: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd3010: dout <= { 2'd1, 8'd024, 10'd194 }; 
        'd3011: dout <= { 2'd2, 8'd010, 10'd344 }; 
        'd3012: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd3013: dout <= { 2'd1, 8'd036, 10'd164 }; 
        'd3014: dout <= { 2'd2, 8'd025, 10'd340 }; 
        'd3015: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd3016: dout <= { 2'd1, 8'd029, 10'd064 }; 
        'd3017: dout <= { 2'd2, 8'd024, 10'd345 }; 
        'd3018: dout <= { 2'd1, 8'd036, 10'd000 }; 
        'd3019: dout <= { 2'd1, 8'd025, 10'd066 }; 
        'd3020: dout <= { 2'd2, 8'd022, 10'd183 }; 
        'd3021: dout <= { 2'd1, 8'd037, 10'd000 }; 
        'd3022: dout <= { 2'd1, 8'd001, 10'd209 }; 
        'd3023: dout <= { 2'd2, 8'd021, 10'd106 }; 
        'd3024: dout <= { 2'd1, 8'd038, 10'd000 }; 
        'd3025: dout <= { 2'd1, 8'd041, 10'd246 }; 
        'd3026: dout <= { 2'd2, 8'd039, 10'd107 }; 
        'd3027: dout <= { 2'd1, 8'd039, 10'd000 }; 
        'd3028: dout <= { 2'd1, 8'd022, 10'd062 }; 
        'd3029: dout <= { 2'd2, 8'd016, 10'd189 }; 
        'd3030: dout <= { 2'd1, 8'd040, 10'd000 }; 
        'd3031: dout <= { 2'd1, 8'd016, 10'd188 }; 
        'd3032: dout <= { 2'd2, 8'd002, 10'd327 }; 
        'd3033: dout <= { 2'd1, 8'd041, 10'd000 }; 
        'd3034: dout <= { 2'd1, 8'd035, 10'd173 }; 
        'd3035: dout <= { 2'd2, 8'd015, 10'd341 }; 
        'd3036: dout <= { 2'd1, 8'd042, 10'd000 }; 
        'd3037: dout <= { 2'd1, 8'd009, 10'd026 }; 
        'd3038: dout <= { 2'd2, 8'd019, 10'd176 }; 
        'd3039: dout <= { 2'd1, 8'd043, 10'd000 }; 
        'd3040: dout <= { 2'd1, 8'd017, 10'd052 }; 
        'd3041: dout <= { 2'd2, 8'd038, 10'd192 }; 
        'd3042: dout <= { 2'd1, 8'd044, 10'd000 }; 
        'd3043: dout <= { 2'd1, 8'd008, 10'd171 }; 
        'd3044: dout <= { 2'd2, 8'd006, 10'd138 }; 
        'd3045: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd3046: dout <= { 2'd1, 8'd012, 10'd077 }; 
        'd3047: dout <= { 2'd2, 8'd002, 10'd157 }; 
        'd3048: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd3049: dout <= { 2'd1, 8'd016, 10'd087 }; 
        'd3050: dout <= { 2'd2, 8'd030, 10'd307 }; 
        'd3051: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd3052: dout <= { 2'd1, 8'd025, 10'd170 }; 
        'd3053: dout <= { 2'd2, 8'd029, 10'd286 }; 
        'd3054: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd3055: dout <= { 2'd1, 8'd044, 10'd038 }; 
        'd3056: dout <= { 2'd2, 8'd042, 10'd181 }; 
        'd3057: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd3058: dout <= { 2'd1, 8'd000, 10'd173 }; 
        'd3059: dout <= { 2'd2, 8'd005, 10'd031 }; 
        'd3060: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd3061: dout <= { 2'd1, 8'd033, 10'd204 }; 
        'd3062: dout <= { 2'd2, 8'd041, 10'd130 }; 
        'd3063: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd3064: dout <= { 2'd1, 8'd019, 10'd055 }; 
        'd3065: dout <= { 2'd2, 8'd008, 10'd171 }; 
        'd3066: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd3067: dout <= { 2'd1, 8'd011, 10'd057 }; 
        'd3068: dout <= { 2'd2, 8'd027, 10'd175 }; 
        'd3069: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd3070: dout <= { 2'd1, 8'd006, 10'd107 }; 
        'd3071: dout <= { 2'd2, 8'd022, 10'd348 }; 
        'd3072: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd3073: dout <= { 2'd1, 8'd031, 10'd231 }; 
        'd3074: dout <= { 2'd2, 8'd010, 10'd265 }; 
        'd3075: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd3076: dout <= { 2'd1, 8'd010, 10'd040 }; 
        'd3077: dout <= { 2'd2, 8'd004, 10'd020 }; 
        'd3078: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd3079: dout <= { 2'd1, 8'd037, 10'd251 }; 
        'd3080: dout <= { 2'd2, 8'd039, 10'd205 }; 
        'd3081: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd3082: dout <= { 2'd1, 8'd017, 10'd251 }; 
        'd3083: dout <= { 2'd2, 8'd015, 10'd079 }; 
        'd3084: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd3085: dout <= { 2'd1, 8'd021, 10'd331 }; 
        'd3086: dout <= { 2'd2, 8'd040, 10'd058 }; 
        'd3087: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd3088: dout <= { 2'd1, 8'd029, 10'd170 }; 
        'd3089: dout <= { 2'd2, 8'd012, 10'd174 }; 
        'd3090: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd3091: dout <= { 2'd1, 8'd014, 10'd135 }; 
        'd3092: dout <= { 2'd2, 8'd034, 10'd290 }; 
        'd3093: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd3094: dout <= { 2'd1, 8'd023, 10'd087 }; 
        'd3095: dout <= { 2'd2, 8'd006, 10'd061 }; 
        'd3096: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd3097: dout <= { 2'd1, 8'd004, 10'd189 }; 
        'd3098: dout <= { 2'd2, 8'd013, 10'd103 }; 
        'd3099: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd3100: dout <= { 2'd1, 8'd009, 10'd271 }; 
        'd3101: dout <= { 2'd2, 8'd007, 10'd198 }; 
        'd3102: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd3103: dout <= { 2'd1, 8'd034, 10'd127 }; 
        'd3104: dout <= { 2'd2, 8'd023, 10'd276 }; 
        'd3105: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd3106: dout <= { 2'd1, 8'd013, 10'd280 }; 
        'd3107: dout <= { 2'd2, 8'd021, 10'd098 }; 
        'd3108: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd3109: dout <= { 2'd1, 8'd039, 10'd029 }; 
        'd3110: dout <= { 2'd2, 8'd009, 10'd089 }; 
        'd3111: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd3112: dout <= { 2'd1, 8'd028, 10'd188 }; 
        'd3113: dout <= { 2'd2, 8'd035, 10'd307 }; 
        'd3114: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd3115: dout <= { 2'd1, 8'd020, 10'd038 }; 
        'd3116: dout <= { 2'd2, 8'd001, 10'd331 }; 
        'd3117: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd3118: dout <= { 2'd1, 8'd002, 10'd332 }; 
        'd3119: dout <= { 2'd2, 8'd016, 10'd158 }; 
        'd3120: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd3121: dout <= { 2'd1, 8'd043, 10'd332 }; 
        'd3122: dout <= { 2'd2, 8'd043, 10'd196 }; 
        'd3123: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd3124: dout <= { 2'd1, 8'd008, 10'd146 }; 
        'd3125: dout <= { 2'd2, 8'd014, 10'd190 }; 
        'd3126: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd3127: dout <= { 2'd1, 8'd042, 10'd109 }; 
        'd3128: dout <= { 2'd2, 8'd036, 10'd008 }; 
        'd3129: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd3130: dout <= { 2'd1, 8'd027, 10'd006 }; 
        'd3131: dout <= { 2'd2, 8'd025, 10'd284 }; 
        'd3132: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd3133: dout <= { 2'd1, 8'd018, 10'd308 }; 
        'd3134: dout <= { 2'd2, 8'd032, 10'd148 }; 
        'd3135: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd3136: dout <= { 2'd1, 8'd022, 10'd263 }; 
        'd3137: dout <= { 2'd2, 8'd026, 10'd248 }; 
        'd3138: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd3139: dout <= { 2'd1, 8'd040, 10'd319 }; 
        'd3140: dout <= { 2'd2, 8'd018, 10'd255 }; 
        'd3141: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd3142: dout <= { 2'd1, 8'd035, 10'd358 }; 
        'd3143: dout <= { 2'd2, 8'd011, 10'd272 }; 
        'd3144: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd3145: dout <= { 2'd1, 8'd007, 10'd299 }; 
        'd3146: dout <= { 2'd2, 8'd003, 10'd165 }; 
        'd3147: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd3148: dout <= { 2'd1, 8'd036, 10'd322 }; 
        'd3149: dout <= { 2'd2, 8'd024, 10'd291 }; 
        'd3150: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd3151: dout <= { 2'd1, 8'd015, 10'd056 }; 
        'd3152: dout <= { 2'd2, 8'd038, 10'd249 }; 
        'd3153: dout <= { 2'd1, 8'd036, 10'd000 }; 
        'd3154: dout <= { 2'd1, 8'd030, 10'd143 }; 
        'd3155: dout <= { 2'd2, 8'd000, 10'd282 }; 
        'd3156: dout <= { 2'd1, 8'd037, 10'd000 }; 
        'd3157: dout <= { 2'd1, 8'd032, 10'd152 }; 
        'd3158: dout <= { 2'd2, 8'd019, 10'd207 }; 
        'd3159: dout <= { 2'd1, 8'd038, 10'd000 }; 
        'd3160: dout <= { 2'd1, 8'd026, 10'd341 }; 
        'd3161: dout <= { 2'd2, 8'd028, 10'd311 }; 
        'd3162: dout <= { 2'd1, 8'd039, 10'd000 }; 
        'd3163: dout <= { 2'd1, 8'd001, 10'd180 }; 
        'd3164: dout <= { 2'd2, 8'd017, 10'd226 }; 
        'd3165: dout <= { 2'd1, 8'd040, 10'd000 }; 
        'd3166: dout <= { 2'd1, 8'd038, 10'd265 }; 
        'd3167: dout <= { 2'd2, 8'd033, 10'd107 }; 
        'd3168: dout <= { 2'd1, 8'd041, 10'd000 }; 
        'd3169: dout <= { 2'd1, 8'd005, 10'd336 }; 
        'd3170: dout <= { 2'd2, 8'd044, 10'd135 }; 
        'd3171: dout <= { 2'd1, 8'd042, 10'd000 }; 
        'd3172: dout <= { 2'd1, 8'd041, 10'd178 }; 
        'd3173: dout <= { 2'd2, 8'd020, 10'd321 }; 
        'd3174: dout <= { 2'd1, 8'd043, 10'd000 }; 
        'd3175: dout <= { 2'd1, 8'd024, 10'd247 }; 
        'd3176: dout <= { 2'd2, 8'd037, 10'd114 }; 
        'd3177: dout <= { 2'd1, 8'd044, 10'd000 }; 
        'd3178: dout <= { 2'd1, 8'd003, 10'd064 }; 
        'd3179: dout <= { 2'd3, 8'd031, 10'd322 }; 
        // Q=36, BaseAddr=3180
        'd3180: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd3181: dout <= { 2'd1, 8'd005, 10'd004 }; 
        'd3182: dout <= { 2'd1, 8'd016, 10'd311 }; 
        'd3183: dout <= { 2'd1, 8'd031, 10'd154 }; 
        'd3184: dout <= { 2'd1, 8'd024, 10'd176 }; 
        'd3185: dout <= { 2'd1, 8'd031, 10'd348 }; 
        'd3186: dout <= { 2'd1, 8'd008, 10'd225 }; 
        'd3187: dout <= { 2'd1, 8'd009, 10'd236 }; 
        'd3188: dout <= { 2'd1, 8'd012, 10'd011 }; 
        'd3189: dout <= { 2'd1, 8'd018, 10'd278 }; 
        'd3190: dout <= { 2'd2, 8'd012, 10'd356 }; 
        'd3191: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd3192: dout <= { 2'd1, 8'd017, 10'd145 }; 
        'd3193: dout <= { 2'd1, 8'd022, 10'd013 }; 
        'd3194: dout <= { 2'd1, 8'd021, 10'd296 }; 
        'd3195: dout <= { 2'd1, 8'd030, 10'd138 }; 
        'd3196: dout <= { 2'd1, 8'd017, 10'd107 }; 
        'd3197: dout <= { 2'd1, 8'd026, 10'd103 }; 
        'd3198: dout <= { 2'd1, 8'd032, 10'd085 }; 
        'd3199: dout <= { 2'd1, 8'd017, 10'd097 }; 
        'd3200: dout <= { 2'd1, 8'd035, 10'd213 }; 
        'd3201: dout <= { 2'd2, 8'd009, 10'd286 }; 
        'd3202: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd3203: dout <= { 2'd1, 8'd030, 10'd242 }; 
        'd3204: dout <= { 2'd1, 8'd009, 10'd154 }; 
        'd3205: dout <= { 2'd1, 8'd012, 10'd078 }; 
        'd3206: dout <= { 2'd1, 8'd029, 10'd196 }; 
        'd3207: dout <= { 2'd1, 8'd020, 10'd336 }; 
        'd3208: dout <= { 2'd1, 8'd009, 10'd291 }; 
        'd3209: dout <= { 2'd1, 8'd024, 10'd015 }; 
        'd3210: dout <= { 2'd1, 8'd019, 10'd216 }; 
        'd3211: dout <= { 2'd1, 8'd020, 10'd082 }; 
        'd3212: dout <= { 2'd2, 8'd033, 10'd059 }; 
        'd3213: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd3214: dout <= { 2'd1, 8'd035, 10'd074 }; 
        'd3215: dout <= { 2'd1, 8'd020, 10'd119 }; 
        'd3216: dout <= { 2'd1, 8'd034, 10'd231 }; 
        'd3217: dout <= { 2'd1, 8'd028, 10'd019 }; 
        'd3218: dout <= { 2'd1, 8'd033, 10'd078 }; 
        'd3219: dout <= { 2'd1, 8'd010, 10'd090 }; 
        'd3220: dout <= { 2'd1, 8'd015, 10'd131 }; 
        'd3221: dout <= { 2'd1, 8'd025, 10'd280 }; 
        'd3222: dout <= { 2'd1, 8'd013, 10'd014 }; 
        'd3223: dout <= { 2'd2, 8'd028, 10'd208 }; 
        'd3224: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd3225: dout <= { 2'd1, 8'd007, 10'd335 }; 
        'd3226: dout <= { 2'd1, 8'd019, 10'd037 }; 
        'd3227: dout <= { 2'd1, 8'd004, 10'd333 }; 
        'd3228: dout <= { 2'd1, 8'd023, 10'd338 }; 
        'd3229: dout <= { 2'd1, 8'd035, 10'd312 }; 
        'd3230: dout <= { 2'd1, 8'd013, 10'd143 }; 
        'd3231: dout <= { 2'd1, 8'd033, 10'd014 }; 
        'd3232: dout <= { 2'd1, 8'd010, 10'd171 }; 
        'd3233: dout <= { 2'd1, 8'd034, 10'd117 }; 
        'd3234: dout <= { 2'd2, 8'd023, 10'd065 }; 
        'd3235: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd3236: dout <= { 2'd1, 8'd024, 10'd189 }; 
        'd3237: dout <= { 2'd1, 8'd015, 10'd197 }; 
        'd3238: dout <= { 2'd1, 8'd003, 10'd059 }; 
        'd3239: dout <= { 2'd1, 8'd016, 10'd103 }; 
        'd3240: dout <= { 2'd1, 8'd019, 10'd159 }; 
        'd3241: dout <= { 2'd1, 8'd024, 10'd306 }; 
        'd3242: dout <= { 2'd1, 8'd028, 10'd298 }; 
        'd3243: dout <= { 2'd1, 8'd005, 10'd113 }; 
        'd3244: dout <= { 2'd1, 8'd003, 10'd028 }; 
        'd3245: dout <= { 2'd2, 8'd002, 10'd095 }; 
        'd3246: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd3247: dout <= { 2'd1, 8'd027, 10'd312 }; 
        'd3248: dout <= { 2'd1, 8'd028, 10'd033 }; 
        'd3249: dout <= { 2'd1, 8'd022, 10'd264 }; 
        'd3250: dout <= { 2'd1, 8'd026, 10'd040 }; 
        'd3251: dout <= { 2'd1, 8'd016, 10'd300 }; 
        'd3252: dout <= { 2'd1, 8'd004, 10'd026 }; 
        'd3253: dout <= { 2'd1, 8'd000, 10'd104 }; 
        'd3254: dout <= { 2'd1, 8'd007, 10'd078 }; 
        'd3255: dout <= { 2'd1, 8'd022, 10'd319 }; 
        'd3256: dout <= { 2'd2, 8'd017, 10'd321 }; 
        'd3257: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd3258: dout <= { 2'd1, 8'd013, 10'd126 }; 
        'd3259: dout <= { 2'd1, 8'd023, 10'd319 }; 
        'd3260: dout <= { 2'd1, 8'd002, 10'd031 }; 
        'd3261: dout <= { 2'd1, 8'd014, 10'd035 }; 
        'd3262: dout <= { 2'd1, 8'd015, 10'd326 }; 
        'd3263: dout <= { 2'd1, 8'd023, 10'd144 }; 
        'd3264: dout <= { 2'd1, 8'd006, 10'd218 }; 
        'd3265: dout <= { 2'd1, 8'd023, 10'd355 }; 
        'd3266: dout <= { 2'd1, 8'd015, 10'd112 }; 
        'd3267: dout <= { 2'd2, 8'd004, 10'd180 }; 
        'd3268: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd3269: dout <= { 2'd1, 8'd006, 10'd234 }; 
        'd3270: dout <= { 2'd1, 8'd011, 10'd114 }; 
        'd3271: dout <= { 2'd1, 8'd008, 10'd262 }; 
        'd3272: dout <= { 2'd1, 8'd017, 10'd011 }; 
        'd3273: dout <= { 2'd1, 8'd027, 10'd123 }; 
        'd3274: dout <= { 2'd1, 8'd030, 10'd062 }; 
        'd3275: dout <= { 2'd1, 8'd031, 10'd219 }; 
        'd3276: dout <= { 2'd1, 8'd018, 10'd344 }; 
        'd3277: dout <= { 2'd1, 8'd011, 10'd238 }; 
        'd3278: dout <= { 2'd2, 8'd032, 10'd195 }; 
        'd3279: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd3280: dout <= { 2'd1, 8'd033, 10'd107 }; 
        'd3281: dout <= { 2'd1, 8'd018, 10'd253 }; 
        'd3282: dout <= { 2'd1, 8'd013, 10'd157 }; 
        'd3283: dout <= { 2'd1, 8'd005, 10'd125 }; 
        'd3284: dout <= { 2'd1, 8'd003, 10'd065 }; 
        'd3285: dout <= { 2'd1, 8'd001, 10'd007 }; 
        'd3286: dout <= { 2'd1, 8'd027, 10'd130 }; 
        'd3287: dout <= { 2'd1, 8'd034, 10'd103 }; 
        'd3288: dout <= { 2'd1, 8'd026, 10'd115 }; 
        'd3289: dout <= { 2'd2, 8'd008, 10'd043 }; 
        'd3290: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd3291: dout <= { 2'd1, 8'd012, 10'd047 }; 
        'd3292: dout <= { 2'd1, 8'd008, 10'd248 }; 
        'd3293: dout <= { 2'd1, 8'd007, 10'd188 }; 
        'd3294: dout <= { 2'd1, 8'd035, 10'd239 }; 
        'd3295: dout <= { 2'd1, 8'd007, 10'd227 }; 
        'd3296: dout <= { 2'd1, 8'd034, 10'd220 }; 
        'd3297: dout <= { 2'd1, 8'd026, 10'd228 }; 
        'd3298: dout <= { 2'd1, 8'd002, 10'd218 }; 
        'd3299: dout <= { 2'd1, 8'd027, 10'd246 }; 
        'd3300: dout <= { 2'd2, 8'd001, 10'd242 }; 
        'd3301: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd3302: dout <= { 2'd1, 8'd016, 10'd325 }; 
        'd3303: dout <= { 2'd1, 8'd024, 10'd120 }; 
        'd3304: dout <= { 2'd1, 8'd015, 10'd252 }; 
        'd3305: dout <= { 2'd1, 8'd032, 10'd312 }; 
        'd3306: dout <= { 2'd1, 8'd006, 10'd063 }; 
        'd3307: dout <= { 2'd1, 8'd012, 10'd245 }; 
        'd3308: dout <= { 2'd1, 8'd003, 10'd254 }; 
        'd3309: dout <= { 2'd1, 8'd014, 10'd331 }; 
        'd3310: dout <= { 2'd1, 8'd006, 10'd168 }; 
        'd3311: dout <= { 2'd2, 8'd019, 10'd151 }; 
        'd3312: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd3313: dout <= { 2'd1, 8'd015, 10'd203 }; 
        'd3314: dout <= { 2'd1, 8'd010, 10'd110 }; 
        'd3315: dout <= { 2'd1, 8'd033, 10'd286 }; 
        'd3316: dout <= { 2'd1, 8'd010, 10'd060 }; 
        'd3317: dout <= { 2'd1, 8'd018, 10'd229 }; 
        'd3318: dout <= { 2'd1, 8'd002, 10'd107 }; 
        'd3319: dout <= { 2'd1, 8'd035, 10'd057 }; 
        'd3320: dout <= { 2'd1, 8'd011, 10'd358 }; 
        'd3321: dout <= { 2'd1, 8'd029, 10'd263 }; 
        'd3322: dout <= { 2'd2, 8'd000, 10'd325 }; 
        'd3323: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd3324: dout <= { 2'd1, 8'd026, 10'd122 }; 
        'd3325: dout <= { 2'd1, 8'd027, 10'd040 }; 
        'd3326: dout <= { 2'd1, 8'd006, 10'd069 }; 
        'd3327: dout <= { 2'd1, 8'd009, 10'd162 }; 
        'd3328: dout <= { 2'd1, 8'd025, 10'd022 }; 
        'd3329: dout <= { 2'd1, 8'd005, 10'd318 }; 
        'd3330: dout <= { 2'd1, 8'd029, 10'd014 }; 
        'd3331: dout <= { 2'd1, 8'd021, 10'd311 }; 
        'd3332: dout <= { 2'd1, 8'd010, 10'd332 }; 
        'd3333: dout <= { 2'd2, 8'd031, 10'd145 }; 
        'd3334: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd3335: dout <= { 2'd1, 8'd029, 10'd042 }; 
        'd3336: dout <= { 2'd1, 8'd025, 10'd125 }; 
        'd3337: dout <= { 2'd1, 8'd020, 10'd221 }; 
        'd3338: dout <= { 2'd1, 8'd001, 10'd096 }; 
        'd3339: dout <= { 2'd1, 8'd032, 10'd264 }; 
        'd3340: dout <= { 2'd1, 8'd021, 10'd214 }; 
        'd3341: dout <= { 2'd1, 8'd008, 10'd105 }; 
        'd3342: dout <= { 2'd1, 8'd030, 10'd082 }; 
        'd3343: dout <= { 2'd1, 8'd007, 10'd175 }; 
        'd3344: dout <= { 2'd2, 8'd021, 10'd166 }; 
        'd3345: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd3346: dout <= { 2'd1, 8'd000, 10'd319 }; 
        'd3347: dout <= { 2'd1, 8'd003, 10'd076 }; 
        'd3348: dout <= { 2'd1, 8'd027, 10'd111 }; 
        'd3349: dout <= { 2'd1, 8'd011, 10'd336 }; 
        'd3350: dout <= { 2'd1, 8'd000, 10'd181 }; 
        'd3351: dout <= { 2'd1, 8'd011, 10'd015 }; 
        'd3352: dout <= { 2'd1, 8'd016, 10'd071 }; 
        'd3353: dout <= { 2'd1, 8'd004, 10'd184 }; 
        'd3354: dout <= { 2'd1, 8'd014, 10'd226 }; 
        'd3355: dout <= { 2'd2, 8'd024, 10'd273 }; 
        'd3356: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd3357: dout <= { 2'd1, 8'd022, 10'd168 }; 
        'd3358: dout <= { 2'd1, 8'd033, 10'd048 }; 
        'd3359: dout <= { 2'd1, 8'd019, 10'd128 }; 
        'd3360: dout <= { 2'd1, 8'd018, 10'd181 }; 
        'd3361: dout <= { 2'd1, 8'd029, 10'd219 }; 
        'd3362: dout <= { 2'd1, 8'd022, 10'd103 }; 
        'd3363: dout <= { 2'd1, 8'd022, 10'd329 }; 
        'd3364: dout <= { 2'd1, 8'd013, 10'd050 }; 
        'd3365: dout <= { 2'd1, 8'd030, 10'd341 }; 
        'd3366: dout <= { 2'd2, 8'd005, 10'd229 }; 
        'd3367: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd3368: dout <= { 2'd1, 8'd021, 10'd345 }; 
        'd3369: dout <= { 2'd1, 8'd017, 10'd152 }; 
        'd3370: dout <= { 2'd1, 8'd000, 10'd243 }; 
        'd3371: dout <= { 2'd1, 8'd025, 10'd217 }; 
        'd3372: dout <= { 2'd1, 8'd028, 10'd212 }; 
        'd3373: dout <= { 2'd1, 8'd014, 10'd058 }; 
        'd3374: dout <= { 2'd1, 8'd001, 10'd315 }; 
        'd3375: dout <= { 2'd1, 8'd020, 10'd081 }; 
        'd3376: dout <= { 2'd1, 8'd016, 10'd186 }; 
        'd3377: dout <= { 2'd2, 8'd025, 10'd332 }; 
        'd3378: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd3379: dout <= { 2'd1, 8'd003, 10'd282 }; 
        'd3380: dout <= { 2'd2, 8'd034, 10'd116 }; 
        'd3381: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd3382: dout <= { 2'd1, 8'd002, 10'd028 }; 
        'd3383: dout <= { 2'd2, 8'd007, 10'd291 }; 
        'd3384: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd3385: dout <= { 2'd1, 8'd008, 10'd247 }; 
        'd3386: dout <= { 2'd2, 8'd026, 10'd284 }; 
        'd3387: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd3388: dout <= { 2'd1, 8'd019, 10'd284 }; 
        'd3389: dout <= { 2'd2, 8'd002, 10'd341 }; 
        'd3390: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd3391: dout <= { 2'd1, 8'd014, 10'd196 }; 
        'd3392: dout <= { 2'd2, 8'd005, 10'd122 }; 
        'd3393: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd3394: dout <= { 2'd1, 8'd031, 10'd340 }; 
        'd3395: dout <= { 2'd2, 8'd035, 10'd107 }; 
        'd3396: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd3397: dout <= { 2'd1, 8'd028, 10'd332 }; 
        'd3398: dout <= { 2'd2, 8'd032, 10'd189 }; 
        'd3399: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd3400: dout <= { 2'd1, 8'd010, 10'd264 }; 
        'd3401: dout <= { 2'd2, 8'd000, 10'd121 }; 
        'd3402: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd3403: dout <= { 2'd1, 8'd009, 10'd198 }; 
        'd3404: dout <= { 2'd2, 8'd021, 10'd285 }; 
        'd3405: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd3406: dout <= { 2'd1, 8'd001, 10'd330 }; 
        'd3407: dout <= { 2'd2, 8'd006, 10'd070 }; 
        'd3408: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd3409: dout <= { 2'd1, 8'd025, 10'd054 }; 
        'd3410: dout <= { 2'd2, 8'd029, 10'd318 }; 
        'd3411: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd3412: dout <= { 2'd1, 8'd020, 10'd084 }; 
        'd3413: dout <= { 2'd2, 8'd013, 10'd303 }; 
        'd3414: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd3415: dout <= { 2'd1, 8'd004, 10'd062 }; 
        'd3416: dout <= { 2'd2, 8'd012, 10'd242 }; 
        'd3417: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd3418: dout <= { 2'd1, 8'd032, 10'd252 }; 
        'd3419: dout <= { 2'd2, 8'd004, 10'd176 }; 
        'd3420: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd3421: dout <= { 2'd1, 8'd034, 10'd203 }; 
        'd3422: dout <= { 2'd2, 8'd014, 10'd238 }; 
        'd3423: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd3424: dout <= { 2'd1, 8'd011, 10'd324 }; 
        'd3425: dout <= { 2'd2, 8'd001, 10'd289 }; 
        'd3426: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd3427: dout <= { 2'd1, 8'd023, 10'd179 }; 
        'd3428: dout <= { 2'd2, 8'd031, 10'd354 }; 
        'd3429: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd3430: dout <= { 2'd1, 8'd018, 10'd088 }; 
        'd3431: dout <= { 2'd2, 8'd030, 10'd338 }; 
        'd3432: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd3433: dout <= { 2'd1, 8'd009, 10'd267 }; 
        'd3434: dout <= { 2'd2, 8'd033, 10'd317 }; 
        'd3435: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd3436: dout <= { 2'd1, 8'd034, 10'd207 }; 
        'd3437: dout <= { 2'd2, 8'd031, 10'd155 }; 
        'd3438: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd3439: dout <= { 2'd1, 8'd035, 10'd119 }; 
        'd3440: dout <= { 2'd2, 8'd019, 10'd135 }; 
        'd3441: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd3442: dout <= { 2'd1, 8'd000, 10'd061 }; 
        'd3443: dout <= { 2'd2, 8'd020, 10'd009 }; 
        'd3444: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd3445: dout <= { 2'd1, 8'd003, 10'd209 }; 
        'd3446: dout <= { 2'd2, 8'd026, 10'd184 }; 
        'd3447: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd3448: dout <= { 2'd1, 8'd001, 10'd297 }; 
        'd3449: dout <= { 2'd2, 8'd028, 10'd067 }; 
        'd3450: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd3451: dout <= { 2'd1, 8'd023, 10'd187 }; 
        'd3452: dout <= { 2'd2, 8'd006, 10'd075 }; 
        'd3453: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd3454: dout <= { 2'd1, 8'd032, 10'd142 }; 
        'd3455: dout <= { 2'd2, 8'd022, 10'd166 }; 
        'd3456: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd3457: dout <= { 2'd1, 8'd027, 10'd306 }; 
        'd3458: dout <= { 2'd2, 8'd005, 10'd223 }; 
        'd3459: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd3460: dout <= { 2'd1, 8'd022, 10'd134 }; 
        'd3461: dout <= { 2'd2, 8'd007, 10'd123 }; 
        'd3462: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd3463: dout <= { 2'd1, 8'd017, 10'd115 }; 
        'd3464: dout <= { 2'd2, 8'd012, 10'd256 }; 
        'd3465: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd3466: dout <= { 2'd1, 8'd030, 10'd340 }; 
        'd3467: dout <= { 2'd2, 8'd010, 10'd182 }; 
        'd3468: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd3469: dout <= { 2'd1, 8'd002, 10'd332 }; 
        'd3470: dout <= { 2'd2, 8'd032, 10'd210 }; 
        'd3471: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd3472: dout <= { 2'd1, 8'd004, 10'd206 }; 
        'd3473: dout <= { 2'd2, 8'd000, 10'd072 }; 
        'd3474: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd3475: dout <= { 2'd1, 8'd026, 10'd244 }; 
        'd3476: dout <= { 2'd2, 8'd024, 10'd267 }; 
        'd3477: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd3478: dout <= { 2'd1, 8'd005, 10'd019 }; 
        'd3479: dout <= { 2'd2, 8'd030, 10'd150 }; 
        'd3480: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd3481: dout <= { 2'd1, 8'd020, 10'd025 }; 
        'd3482: dout <= { 2'd2, 8'd008, 10'd036 }; 
        'd3483: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd3484: dout <= { 2'd1, 8'd029, 10'd034 }; 
        'd3485: dout <= { 2'd2, 8'd018, 10'd331 }; 
        'd3486: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd3487: dout <= { 2'd1, 8'd019, 10'd265 }; 
        'd3488: dout <= { 2'd2, 8'd004, 10'd167 }; 
        'd3489: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd3490: dout <= { 2'd1, 8'd024, 10'd008 }; 
        'd3491: dout <= { 2'd2, 8'd029, 10'd210 }; 
        'd3492: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd3493: dout <= { 2'd1, 8'd011, 10'd123 }; 
        'd3494: dout <= { 2'd2, 8'd021, 10'd116 }; 
        'd3495: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd3496: dout <= { 2'd1, 8'd006, 10'd111 }; 
        'd3497: dout <= { 2'd2, 8'd015, 10'd265 }; 
        'd3498: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd3499: dout <= { 2'd1, 8'd028, 10'd339 }; 
        'd3500: dout <= { 2'd2, 8'd003, 10'd216 }; 
        'd3501: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd3502: dout <= { 2'd1, 8'd018, 10'd041 }; 
        'd3503: dout <= { 2'd2, 8'd034, 10'd243 }; 
        'd3504: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd3505: dout <= { 2'd1, 8'd021, 10'd298 }; 
        'd3506: dout <= { 2'd2, 8'd009, 10'd110 }; 
        'd3507: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd3508: dout <= { 2'd1, 8'd012, 10'd121 }; 
        'd3509: dout <= { 2'd2, 8'd023, 10'd096 }; 
        'd3510: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd3511: dout <= { 2'd1, 8'd016, 10'd175 }; 
        'd3512: dout <= { 2'd2, 8'd014, 10'd148 }; 
        'd3513: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd3514: dout <= { 2'd1, 8'd007, 10'd068 }; 
        'd3515: dout <= { 2'd2, 8'd001, 10'd097 }; 
        'd3516: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd3517: dout <= { 2'd1, 8'd025, 10'd337 }; 
        'd3518: dout <= { 2'd2, 8'd025, 10'd205 }; 
        'd3519: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd3520: dout <= { 2'd1, 8'd010, 10'd183 }; 
        'd3521: dout <= { 2'd2, 8'd011, 10'd319 }; 
        'd3522: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd3523: dout <= { 2'd1, 8'd033, 10'd327 }; 
        'd3524: dout <= { 2'd2, 8'd027, 10'd123 }; 
        'd3525: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd3526: dout <= { 2'd1, 8'd013, 10'd267 }; 
        'd3527: dout <= { 2'd2, 8'd002, 10'd058 }; 
        'd3528: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd3529: dout <= { 2'd1, 8'd015, 10'd131 }; 
        'd3530: dout <= { 2'd2, 8'd017, 10'd064 }; 
        'd3531: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd3532: dout <= { 2'd1, 8'd014, 10'd099 }; 
        'd3533: dout <= { 2'd2, 8'd016, 10'd072 }; 
        'd3534: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd3535: dout <= { 2'd1, 8'd008, 10'd236 }; 
        'd3536: dout <= { 2'd2, 8'd013, 10'd051 }; 
        'd3537: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd3538: dout <= { 2'd1, 8'd031, 10'd111 }; 
        'd3539: dout <= { 2'd2, 8'd035, 10'd031 }; 
        'd3540: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd3541: dout <= { 2'd1, 8'd031, 10'd156 }; 
        'd3542: dout <= { 2'd2, 8'd003, 10'd137 }; 
        'd3543: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd3544: dout <= { 2'd1, 8'd007, 10'd117 }; 
        'd3545: dout <= { 2'd2, 8'd034, 10'd051 }; 
        'd3546: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd3547: dout <= { 2'd1, 8'd024, 10'd304 }; 
        'd3548: dout <= { 2'd2, 8'd026, 10'd223 }; 
        'd3549: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd3550: dout <= { 2'd1, 8'd022, 10'd193 }; 
        'd3551: dout <= { 2'd2, 8'd011, 10'd151 }; 
        'd3552: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd3553: dout <= { 2'd1, 8'd013, 10'd089 }; 
        'd3554: dout <= { 2'd2, 8'd022, 10'd156 }; 
        'd3555: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd3556: dout <= { 2'd1, 8'd008, 10'd249 }; 
        'd3557: dout <= { 2'd2, 8'd021, 10'd018 }; 
        'd3558: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd3559: dout <= { 2'd1, 8'd002, 10'd156 }; 
        'd3560: dout <= { 2'd2, 8'd016, 10'd346 }; 
        'd3561: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd3562: dout <= { 2'd1, 8'd017, 10'd040 }; 
        'd3563: dout <= { 2'd2, 8'd020, 10'd035 }; 
        'd3564: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd3565: dout <= { 2'd1, 8'd012, 10'd246 }; 
        'd3566: dout <= { 2'd2, 8'd031, 10'd107 }; 
        'd3567: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd3568: dout <= { 2'd1, 8'd010, 10'd246 }; 
        'd3569: dout <= { 2'd2, 8'd000, 10'd034 }; 
        'd3570: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd3571: dout <= { 2'd1, 8'd019, 10'd232 }; 
        'd3572: dout <= { 2'd2, 8'd032, 10'd165 }; 
        'd3573: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd3574: dout <= { 2'd1, 8'd014, 10'd007 }; 
        'd3575: dout <= { 2'd2, 8'd013, 10'd122 }; 
        'd3576: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd3577: dout <= { 2'd1, 8'd034, 10'd102 }; 
        'd3578: dout <= { 2'd2, 8'd004, 10'd090 }; 
        'd3579: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd3580: dout <= { 2'd1, 8'd027, 10'd167 }; 
        'd3581: dout <= { 2'd2, 8'd012, 10'd162 }; 
        'd3582: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd3583: dout <= { 2'd1, 8'd000, 10'd200 }; 
        'd3584: dout <= { 2'd2, 8'd007, 10'd091 }; 
        'd3585: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd3586: dout <= { 2'd1, 8'd026, 10'd041 }; 
        'd3587: dout <= { 2'd2, 8'd014, 10'd313 }; 
        'd3588: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd3589: dout <= { 2'd1, 8'd006, 10'd342 }; 
        'd3590: dout <= { 2'd2, 8'd006, 10'd061 }; 
        'd3591: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd3592: dout <= { 2'd1, 8'd023, 10'd125 }; 
        'd3593: dout <= { 2'd2, 8'd029, 10'd026 }; 
        'd3594: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd3595: dout <= { 2'd1, 8'd011, 10'd266 }; 
        'd3596: dout <= { 2'd2, 8'd027, 10'd194 }; 
        'd3597: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd3598: dout <= { 2'd1, 8'd032, 10'd070 }; 
        'd3599: dout <= { 2'd2, 8'd035, 10'd056 }; 
        'd3600: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd3601: dout <= { 2'd1, 8'd021, 10'd334 }; 
        'd3602: dout <= { 2'd2, 8'd010, 10'd286 }; 
        'd3603: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd3604: dout <= { 2'd1, 8'd018, 10'd307 }; 
        'd3605: dout <= { 2'd2, 8'd028, 10'd141 }; 
        'd3606: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd3607: dout <= { 2'd1, 8'd003, 10'd184 }; 
        'd3608: dout <= { 2'd2, 8'd030, 10'd191 }; 
        'd3609: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd3610: dout <= { 2'd1, 8'd025, 10'd274 }; 
        'd3611: dout <= { 2'd2, 8'd033, 10'd058 }; 
        'd3612: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd3613: dout <= { 2'd1, 8'd001, 10'd023 }; 
        'd3614: dout <= { 2'd2, 8'd017, 10'd269 }; 
        'd3615: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd3616: dout <= { 2'd1, 8'd005, 10'd061 }; 
        'd3617: dout <= { 2'd2, 8'd019, 10'd050 }; 
        'd3618: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd3619: dout <= { 2'd1, 8'd029, 10'd185 }; 
        'd3620: dout <= { 2'd2, 8'd001, 10'd359 }; 
        'd3621: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd3622: dout <= { 2'd1, 8'd015, 10'd059 }; 
        'd3623: dout <= { 2'd2, 8'd009, 10'd243 }; 
        'd3624: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd3625: dout <= { 2'd1, 8'd016, 10'd333 }; 
        'd3626: dout <= { 2'd2, 8'd008, 10'd165 }; 
        'd3627: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd3628: dout <= { 2'd1, 8'd028, 10'd241 }; 
        'd3629: dout <= { 2'd2, 8'd023, 10'd088 }; 
        'd3630: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd3631: dout <= { 2'd1, 8'd035, 10'd226 }; 
        'd3632: dout <= { 2'd2, 8'd025, 10'd303 }; 
        'd3633: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd3634: dout <= { 2'd1, 8'd033, 10'd174 }; 
        'd3635: dout <= { 2'd2, 8'd024, 10'd197 }; 
        'd3636: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd3637: dout <= { 2'd1, 8'd004, 10'd017 }; 
        'd3638: dout <= { 2'd2, 8'd018, 10'd198 }; 
        'd3639: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd3640: dout <= { 2'd1, 8'd030, 10'd142 }; 
        'd3641: dout <= { 2'd2, 8'd005, 10'd271 }; 
        'd3642: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd3643: dout <= { 2'd1, 8'd009, 10'd288 }; 
        'd3644: dout <= { 2'd2, 8'd002, 10'd226 }; 
        'd3645: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd3646: dout <= { 2'd1, 8'd020, 10'd211 }; 
        'd3647: dout <= { 2'd2, 8'd015, 10'd161 }; 
        'd3648: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd3649: dout <= { 2'd1, 8'd013, 10'd202 }; 
        'd3650: dout <= { 2'd2, 8'd035, 10'd273 }; 
        'd3651: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd3652: dout <= { 2'd1, 8'd024, 10'd215 }; 
        'd3653: dout <= { 2'd2, 8'd031, 10'd301 }; 
        'd3654: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd3655: dout <= { 2'd1, 8'd031, 10'd342 }; 
        'd3656: dout <= { 2'd2, 8'd019, 10'd250 }; 
        'd3657: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd3658: dout <= { 2'd1, 8'd022, 10'd122 }; 
        'd3659: dout <= { 2'd2, 8'd015, 10'd231 }; 
        'd3660: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd3661: dout <= { 2'd1, 8'd008, 10'd096 }; 
        'd3662: dout <= { 2'd2, 8'd030, 10'd017 }; 
        'd3663: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd3664: dout <= { 2'd1, 8'd012, 10'd193 }; 
        'd3665: dout <= { 2'd2, 8'd023, 10'd056 }; 
        'd3666: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd3667: dout <= { 2'd1, 8'd030, 10'd021 }; 
        'd3668: dout <= { 2'd2, 8'd033, 10'd083 }; 
        'd3669: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd3670: dout <= { 2'd1, 8'd026, 10'd019 }; 
        'd3671: dout <= { 2'd2, 8'd034, 10'd057 }; 
        'd3672: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd3673: dout <= { 2'd1, 8'd007, 10'd206 }; 
        'd3674: dout <= { 2'd2, 8'd021, 10'd155 }; 
        'd3675: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd3676: dout <= { 2'd1, 8'd020, 10'd225 }; 
        'd3677: dout <= { 2'd2, 8'd025, 10'd135 }; 
        'd3678: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd3679: dout <= { 2'd1, 8'd001, 10'd344 }; 
        'd3680: dout <= { 2'd2, 8'd002, 10'd333 }; 
        'd3681: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd3682: dout <= { 2'd1, 8'd019, 10'd270 }; 
        'd3683: dout <= { 2'd2, 8'd026, 10'd278 }; 
        'd3684: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd3685: dout <= { 2'd1, 8'd028, 10'd011 }; 
        'd3686: dout <= { 2'd2, 8'd010, 10'd282 }; 
        'd3687: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd3688: dout <= { 2'd1, 8'd015, 10'd037 }; 
        'd3689: dout <= { 2'd2, 8'd001, 10'd211 }; 
        'd3690: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd3691: dout <= { 2'd1, 8'd010, 10'd040 }; 
        'd3692: dout <= { 2'd2, 8'd004, 10'd003 }; 
        'd3693: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd3694: dout <= { 2'd1, 8'd009, 10'd221 }; 
        'd3695: dout <= { 2'd2, 8'd018, 10'd235 }; 
        'd3696: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd3697: dout <= { 2'd1, 8'd017, 10'd248 }; 
        'd3698: dout <= { 2'd2, 8'd017, 10'd205 }; 
        'd3699: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd3700: dout <= { 2'd1, 8'd002, 10'd183 }; 
        'd3701: dout <= { 2'd2, 8'd000, 10'd231 }; 
        'd3702: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd3703: dout <= { 2'd1, 8'd034, 10'd189 }; 
        'd3704: dout <= { 2'd2, 8'd011, 10'd250 }; 
        'd3705: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd3706: dout <= { 2'd1, 8'd018, 10'd171 }; 
        'd3707: dout <= { 2'd2, 8'd014, 10'd261 }; 
        'd3708: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd3709: dout <= { 2'd1, 8'd003, 10'd007 }; 
        'd3710: dout <= { 2'd2, 8'd005, 10'd003 }; 
        'd3711: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd3712: dout <= { 2'd1, 8'd005, 10'd172 }; 
        'd3713: dout <= { 2'd2, 8'd003, 10'd162 }; 
        'd3714: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd3715: dout <= { 2'd1, 8'd014, 10'd358 }; 
        'd3716: dout <= { 2'd2, 8'd028, 10'd106 }; 
        'd3717: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd3718: dout <= { 2'd1, 8'd021, 10'd121 }; 
        'd3719: dout <= { 2'd2, 8'd013, 10'd097 }; 
        'd3720: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd3721: dout <= { 2'd1, 8'd006, 10'd152 }; 
        'd3722: dout <= { 2'd2, 8'd032, 10'd240 }; 
        'd3723: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd3724: dout <= { 2'd1, 8'd025, 10'd123 }; 
        'd3725: dout <= { 2'd2, 8'd008, 10'd059 }; 
        'd3726: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd3727: dout <= { 2'd1, 8'd004, 10'd270 }; 
        'd3728: dout <= { 2'd2, 8'd012, 10'd038 }; 
        'd3729: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd3730: dout <= { 2'd1, 8'd035, 10'd336 }; 
        'd3731: dout <= { 2'd2, 8'd006, 10'd320 }; 
        'd3732: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd3733: dout <= { 2'd1, 8'd011, 10'd342 }; 
        'd3734: dout <= { 2'd2, 8'd007, 10'd264 }; 
        'd3735: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd3736: dout <= { 2'd1, 8'd023, 10'd228 }; 
        'd3737: dout <= { 2'd2, 8'd024, 10'd048 }; 
        'd3738: dout <= { 2'd1, 8'd030, 10'd000 }; 
        'd3739: dout <= { 2'd1, 8'd029, 10'd013 }; 
        'd3740: dout <= { 2'd2, 8'd022, 10'd250 }; 
        'd3741: dout <= { 2'd1, 8'd031, 10'd000 }; 
        'd3742: dout <= { 2'd1, 8'd000, 10'd258 }; 
        'd3743: dout <= { 2'd2, 8'd020, 10'd085 }; 
        'd3744: dout <= { 2'd1, 8'd032, 10'd000 }; 
        'd3745: dout <= { 2'd1, 8'd033, 10'd068 }; 
        'd3746: dout <= { 2'd2, 8'd027, 10'd208 }; 
        'd3747: dout <= { 2'd1, 8'd033, 10'd000 }; 
        'd3748: dout <= { 2'd1, 8'd032, 10'd074 }; 
        'd3749: dout <= { 2'd2, 8'd016, 10'd007 }; 
        'd3750: dout <= { 2'd1, 8'd034, 10'd000 }; 
        'd3751: dout <= { 2'd1, 8'd027, 10'd111 }; 
        'd3752: dout <= { 2'd2, 8'd029, 10'd342 }; 
        'd3753: dout <= { 2'd1, 8'd035, 10'd000 }; 
        'd3754: dout <= { 2'd1, 8'd016, 10'd197 }; 
        'd3755: dout <= { 2'd3, 8'd009, 10'd154 }; 
        // Q=30, BaseAddr=3756
        'd3756: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd3757: dout <= { 2'd1, 8'd012, 10'd145 }; 
        'd3758: dout <= { 2'd1, 8'd026, 10'd013 }; 
        'd3759: dout <= { 2'd1, 8'd029, 10'd296 }; 
        'd3760: dout <= { 2'd1, 8'd016, 10'd138 }; 
        'd3761: dout <= { 2'd1, 8'd006, 10'd107 }; 
        'd3762: dout <= { 2'd1, 8'd022, 10'd103 }; 
        'd3763: dout <= { 2'd1, 8'd010, 10'd085 }; 
        'd3764: dout <= { 2'd1, 8'd002, 10'd097 }; 
        'd3765: dout <= { 2'd1, 8'd015, 10'd213 }; 
        'd3766: dout <= { 2'd1, 8'd013, 10'd286 }; 
        'd3767: dout <= { 2'd1, 8'd019, 10'd165 }; 
        'd3768: dout <= { 2'd2, 8'd003, 10'd224 }; 
        'd3769: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd3770: dout <= { 2'd1, 8'd019, 10'd082 }; 
        'd3771: dout <= { 2'd1, 8'd016, 10'd059 }; 
        'd3772: dout <= { 2'd1, 8'd008, 10'd299 }; 
        'd3773: dout <= { 2'd1, 8'd011, 10'd100 }; 
        'd3774: dout <= { 2'd1, 8'd019, 10'd144 }; 
        'd3775: dout <= { 2'd1, 8'd013, 10'd310 }; 
        'd3776: dout <= { 2'd1, 8'd007, 10'd213 }; 
        'd3777: dout <= { 2'd1, 8'd017, 10'd098 }; 
        'd3778: dout <= { 2'd1, 8'd028, 10'd242 }; 
        'd3779: dout <= { 2'd1, 8'd024, 10'd182 }; 
        'd3780: dout <= { 2'd1, 8'd001, 10'd201 }; 
        'd3781: dout <= { 2'd2, 8'd017, 10'd340 }; 
        'd3782: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd3783: dout <= { 2'd1, 8'd005, 10'd339 }; 
        'd3784: dout <= { 2'd1, 8'd009, 10'd300 }; 
        'd3785: dout <= { 2'd1, 8'd019, 10'd329 }; 
        'd3786: dout <= { 2'd1, 8'd001, 10'd103 }; 
        'd3787: dout <= { 2'd1, 8'd005, 10'd166 }; 
        'd3788: dout <= { 2'd1, 8'd007, 10'd242 }; 
        'd3789: dout <= { 2'd1, 8'd012, 10'd136 }; 
        'd3790: dout <= { 2'd1, 8'd024, 10'd295 }; 
        'd3791: dout <= { 2'd1, 8'd001, 10'd189 }; 
        'd3792: dout <= { 2'd1, 8'd017, 10'd092 }; 
        'd3793: dout <= { 2'd1, 8'd029, 10'd072 }; 
        'd3794: dout <= { 2'd2, 8'd016, 10'd290 }; 
        'd3795: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd3796: dout <= { 2'd1, 8'd022, 10'd301 }; 
        'd3797: dout <= { 2'd1, 8'd025, 10'd159 }; 
        'd3798: dout <= { 2'd1, 8'd024, 10'd130 }; 
        'd3799: dout <= { 2'd1, 8'd010, 10'd112 }; 
        'd3800: dout <= { 2'd1, 8'd008, 10'd335 }; 
        'd3801: dout <= { 2'd1, 8'd018, 10'd037 }; 
        'd3802: dout <= { 2'd1, 8'd006, 10'd333 }; 
        'd3803: dout <= { 2'd1, 8'd025, 10'd338 }; 
        'd3804: dout <= { 2'd1, 8'd000, 10'd312 }; 
        'd3805: dout <= { 2'd1, 8'd007, 10'd143 }; 
        'd3806: dout <= { 2'd1, 8'd014, 10'd014 }; 
        'd3807: dout <= { 2'd2, 8'd008, 10'd171 }; 
        'd3808: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd3809: dout <= { 2'd1, 8'd009, 10'd079 }; 
        'd3810: dout <= { 2'd1, 8'd004, 10'd261 }; 
        'd3811: dout <= { 2'd1, 8'd005, 10'd161 }; 
        'd3812: dout <= { 2'd1, 8'd017, 10'd077 }; 
        'd3813: dout <= { 2'd1, 8'd003, 10'd328 }; 
        'd3814: dout <= { 2'd1, 8'd024, 10'd026 }; 
        'd3815: dout <= { 2'd1, 8'd029, 10'd010 }; 
        'd3816: dout <= { 2'd1, 8'd013, 10'd278 }; 
        'd3817: dout <= { 2'd1, 8'd027, 10'd238 }; 
        'd3818: dout <= { 2'd1, 8'd010, 10'd102 }; 
        'd3819: dout <= { 2'd1, 8'd028, 10'd050 }; 
        'd3820: dout <= { 2'd2, 8'd021, 10'd243 }; 
        'd3821: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd3822: dout <= { 2'd1, 8'd015, 10'd114 }; 
        'd3823: dout <= { 2'd1, 8'd011, 10'd262 }; 
        'd3824: dout <= { 2'd1, 8'd018, 10'd011 }; 
        'd3825: dout <= { 2'd1, 8'd003, 10'd123 }; 
        'd3826: dout <= { 2'd1, 8'd016, 10'd062 }; 
        'd3827: dout <= { 2'd1, 8'd015, 10'd219 }; 
        'd3828: dout <= { 2'd1, 8'd020, 10'd344 }; 
        'd3829: dout <= { 2'd1, 8'd004, 10'd238 }; 
        'd3830: dout <= { 2'd1, 8'd020, 10'd195 }; 
        'd3831: dout <= { 2'd1, 8'd014, 10'd069 }; 
        'd3832: dout <= { 2'd1, 8'd002, 10'd135 }; 
        'd3833: dout <= { 2'd2, 8'd020, 10'd092 }; 
        'd3834: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd3835: dout <= { 2'd1, 8'd017, 10'd130 }; 
        'd3836: dout <= { 2'd1, 8'd021, 10'd103 }; 
        'd3837: dout <= { 2'd1, 8'd026, 10'd115 }; 
        'd3838: dout <= { 2'd1, 8'd014, 10'd043 }; 
        'd3839: dout <= { 2'd1, 8'd011, 10'd344 }; 
        'd3840: dout <= { 2'd1, 8'd029, 10'd197 }; 
        'd3841: dout <= { 2'd1, 8'd009, 10'd173 }; 
        'd3842: dout <= { 2'd1, 8'd021, 10'd053 }; 
        'd3843: dout <= { 2'd1, 8'd011, 10'd066 }; 
        'd3844: dout <= { 2'd1, 8'd009, 10'd023 }; 
        'd3845: dout <= { 2'd1, 8'd006, 10'd277 }; 
        'd3846: dout <= { 2'd2, 8'd000, 10'd332 }; 
        'd3847: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd3848: dout <= { 2'd1, 8'd013, 10'd229 }; 
        'd3849: dout <= { 2'd1, 8'd027, 10'd107 }; 
        'd3850: dout <= { 2'd1, 8'd007, 10'd057 }; 
        'd3851: dout <= { 2'd1, 8'd012, 10'd358 }; 
        'd3852: dout <= { 2'd1, 8'd001, 10'd263 }; 
        'd3853: dout <= { 2'd1, 8'd014, 10'd325 }; 
        'd3854: dout <= { 2'd1, 8'd005, 10'd158 }; 
        'd3855: dout <= { 2'd1, 8'd018, 10'd129 }; 
        'd3856: dout <= { 2'd1, 8'd019, 10'd333 }; 
        'd3857: dout <= { 2'd1, 8'd006, 10'd139 }; 
        'd3858: dout <= { 2'd1, 8'd024, 10'd153 }; 
        'd3859: dout <= { 2'd2, 8'd007, 10'd052 }; 
        'd3860: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd3861: dout <= { 2'd1, 8'd027, 10'd352 }; 
        'd3862: dout <= { 2'd1, 8'd005, 10'd073 }; 
        'd3863: dout <= { 2'd1, 8'd009, 10'd056 }; 
        'd3864: dout <= { 2'd1, 8'd028, 10'd098 }; 
        'd3865: dout <= { 2'd1, 8'd020, 10'd180 }; 
        'd3866: dout <= { 2'd1, 8'd000, 10'd086 }; 
        'd3867: dout <= { 2'd1, 8'd003, 10'd096 }; 
        'd3868: dout <= { 2'd1, 8'd016, 10'd216 }; 
        'd3869: dout <= { 2'd1, 8'd021, 10'd003 }; 
        'd3870: dout <= { 2'd1, 8'd023, 10'd200 }; 
        'd3871: dout <= { 2'd1, 8'd004, 10'd034 }; 
        'd3872: dout <= { 2'd2, 8'd009, 10'd148 }; 
        'd3873: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd3874: dout <= { 2'd1, 8'd006, 10'd126 }; 
        'd3875: dout <= { 2'd1, 8'd013, 10'd286 }; 
        'd3876: dout <= { 2'd1, 8'd004, 10'd069 }; 
        'd3877: dout <= { 2'd1, 8'd021, 10'd110 }; 
        'd3878: dout <= { 2'd1, 8'd017, 10'd168 }; 
        'd3879: dout <= { 2'd1, 8'd010, 10'd048 }; 
        'd3880: dout <= { 2'd1, 8'd000, 10'd128 }; 
        'd3881: dout <= { 2'd1, 8'd014, 10'd181 }; 
        'd3882: dout <= { 2'd1, 8'd002, 10'd219 }; 
        'd3883: dout <= { 2'd1, 8'd004, 10'd103 }; 
        'd3884: dout <= { 2'd1, 8'd022, 10'd329 }; 
        'd3885: dout <= { 2'd2, 8'd012, 10'd050 }; 
        'd3886: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd3887: dout <= { 2'd1, 8'd028, 10'd284 }; 
        'd3888: dout <= { 2'd1, 8'd018, 10'd061 }; 
        'd3889: dout <= { 2'd1, 8'd022, 10'd345 }; 
        'd3890: dout <= { 2'd1, 8'd025, 10'd152 }; 
        'd3891: dout <= { 2'd1, 8'd023, 10'd243 }; 
        'd3892: dout <= { 2'd1, 8'd026, 10'd217 }; 
        'd3893: dout <= { 2'd1, 8'd019, 10'd212 }; 
        'd3894: dout <= { 2'd1, 8'd026, 10'd058 }; 
        'd3895: dout <= { 2'd1, 8'd012, 10'd315 }; 
        'd3896: dout <= { 2'd1, 8'd026, 10'd081 }; 
        'd3897: dout <= { 2'd1, 8'd026, 10'd186 }; 
        'd3898: dout <= { 2'd2, 8'd015, 10'd332 }; 
        'd3899: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd3900: dout <= { 2'd1, 8'd014, 10'd273 }; 
        'd3901: dout <= { 2'd1, 8'd003, 10'd353 }; 
        'd3902: dout <= { 2'd1, 8'd015, 10'd264 }; 
        'd3903: dout <= { 2'd1, 8'd006, 10'd121 }; 
        'd3904: dout <= { 2'd1, 8'd012, 10'd129 }; 
        'd3905: dout <= { 2'd1, 8'd004, 10'd013 }; 
        'd3906: dout <= { 2'd1, 8'd028, 10'd198 }; 
        'd3907: dout <= { 2'd1, 8'd011, 10'd285 }; 
        'd3908: dout <= { 2'd1, 8'd025, 10'd079 }; 
        'd3909: dout <= { 2'd1, 8'd029, 10'd242 }; 
        'd3910: dout <= { 2'd1, 8'd027, 10'd308 }; 
        'd3911: dout <= { 2'd2, 8'd018, 10'd332 }; 
        'd3912: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd3913: dout <= { 2'd1, 8'd025, 10'd259 }; 
        'd3914: dout <= { 2'd1, 8'd014, 10'd002 }; 
        'd3915: dout <= { 2'd1, 8'd013, 10'd054 }; 
        'd3916: dout <= { 2'd1, 8'd002, 10'd318 }; 
        'd3917: dout <= { 2'd1, 8'd027, 10'd228 }; 
        'd3918: dout <= { 2'd1, 8'd002, 10'd245 }; 
        'd3919: dout <= { 2'd1, 8'd027, 10'd213 }; 
        'd3920: dout <= { 2'd1, 8'd008, 10'd252 }; 
        'd3921: dout <= { 2'd1, 8'd003, 10'd354 }; 
        'd3922: dout <= { 2'd1, 8'd005, 10'd024 }; 
        'd3923: dout <= { 2'd1, 8'd011, 10'd084 }; 
        'd3924: dout <= { 2'd2, 8'd025, 10'd303 }; 
        'd3925: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd3926: dout <= { 2'd1, 8'd011, 10'd238 }; 
        'd3927: dout <= { 2'd1, 8'd022, 10'd082 }; 
        'd3928: dout <= { 2'd1, 8'd000, 10'd142 }; 
        'd3929: dout <= { 2'd1, 8'd023, 10'd166 }; 
        'd3930: dout <= { 2'd1, 8'd025, 10'd336 }; 
        'd3931: dout <= { 2'd1, 8'd009, 10'd247 }; 
        'd3932: dout <= { 2'd1, 8'd023, 10'd306 }; 
        'd3933: dout <= { 2'd1, 8'd001, 10'd223 }; 
        'd3934: dout <= { 2'd1, 8'd008, 10'd293 }; 
        'd3935: dout <= { 2'd1, 8'd022, 10'd069 }; 
        'd3936: dout <= { 2'd1, 8'd013, 10'd275 }; 
        'd3937: dout <= { 2'd2, 8'd005, 10'd125 }; 
        'd3938: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd3939: dout <= { 2'd1, 8'd000, 10'd120 }; 
        'd3940: dout <= { 2'd1, 8'd000, 10'd019 }; 
        'd3941: dout <= { 2'd1, 8'd027, 10'd150 }; 
        'd3942: dout <= { 2'd1, 8'd020, 10'd006 }; 
        'd3943: dout <= { 2'd1, 8'd028, 10'd323 }; 
        'd3944: dout <= { 2'd1, 8'd021, 10'd225 }; 
        'd3945: dout <= { 2'd1, 8'd015, 10'd066 }; 
        'd3946: dout <= { 2'd1, 8'd022, 10'd296 }; 
        'd3947: dout <= { 2'd1, 8'd016, 10'd181 }; 
        'd3948: dout <= { 2'd1, 8'd018, 10'd025 }; 
        'd3949: dout <= { 2'd1, 8'd023, 10'd036 }; 
        'd3950: dout <= { 2'd2, 8'd010, 10'd217 }; 
        'd3951: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd3952: dout <= { 2'd1, 8'd004, 10'd210 }; 
        'd3953: dout <= { 2'd2, 8'd001, 10'd254 }; 
        'd3954: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd3955: dout <= { 2'd1, 8'd018, 10'd216 }; 
        'd3956: dout <= { 2'd2, 8'd029, 10'd306 }; 
        'd3957: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd3958: dout <= { 2'd1, 8'd003, 10'd243 }; 
        'd3959: dout <= { 2'd2, 8'd006, 10'd226 }; 
        'd3960: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd3961: dout <= { 2'd1, 8'd010, 10'd198 }; 
        'd3962: dout <= { 2'd2, 8'd028, 10'd056 }; 
        'd3963: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd3964: dout <= { 2'd1, 8'd001, 10'd284 }; 
        'd3965: dout <= { 2'd2, 8'd023, 10'd059 }; 
        'd3966: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd3967: dout <= { 2'd1, 8'd024, 10'd205 }; 
        'd3968: dout <= { 2'd2, 8'd024, 10'd261 }; 
        'd3969: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd3970: dout <= { 2'd1, 8'd023, 10'd325 }; 
        'd3971: dout <= { 2'd2, 8'd020, 10'd039 }; 
        'd3972: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd3973: dout <= { 2'd1, 8'd007, 10'd317 }; 
        'd3974: dout <= { 2'd2, 8'd008, 10'd342 }; 
        'd3975: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd3976: dout <= { 2'd1, 8'd021, 10'd072 }; 
        'd3977: dout <= { 2'd2, 8'd019, 10'd311 }; 
        'd3978: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd3979: dout <= { 2'd1, 8'd029, 10'd064 }; 
        'd3980: dout <= { 2'd2, 8'd010, 10'd185 }; 
        'd3981: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd3982: dout <= { 2'd1, 8'd026, 10'd051 }; 
        'd3983: dout <= { 2'd2, 8'd015, 10'd018 }; 
        'd3984: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd3985: dout <= { 2'd1, 8'd020, 10'd286 }; 
        'd3986: dout <= { 2'd2, 8'd017, 10'd127 }; 
        'd3987: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd3988: dout <= { 2'd1, 8'd002, 10'd169 }; 
        'd3989: dout <= { 2'd2, 8'd007, 10'd035 }; 
        'd3990: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd3991: dout <= { 2'd1, 8'd008, 10'd264 }; 
        'd3992: dout <= { 2'd2, 8'd002, 10'd118 }; 
        'd3993: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd3994: dout <= { 2'd1, 8'd016, 10'd107 }; 
        'd3995: dout <= { 2'd2, 8'd012, 10'd125 }; 
        'd3996: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd3997: dout <= { 2'd1, 8'd025, 10'd234 }; 
        'd3998: dout <= { 2'd2, 8'd020, 10'd080 }; 
        'd3999: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4000: dout <= { 2'd1, 8'd015, 10'd321 }; 
        'd4001: dout <= { 2'd2, 8'd001, 10'd088 }; 
        'd4002: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4003: dout <= { 2'd1, 8'd014, 10'd092 }; 
        'd4004: dout <= { 2'd2, 8'd022, 10'd081 }; 
        'd4005: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4006: dout <= { 2'd1, 8'd021, 10'd177 }; 
        'd4007: dout <= { 2'd2, 8'd021, 10'd067 }; 
        'd4008: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4009: dout <= { 2'd1, 8'd010, 10'd313 }; 
        'd4010: dout <= { 2'd2, 8'd003, 10'd250 }; 
        'd4011: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4012: dout <= { 2'd1, 8'd020, 10'd061 }; 
        'd4013: dout <= { 2'd2, 8'd028, 10'd077 }; 
        'd4014: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4015: dout <= { 2'd1, 8'd016, 10'd348 }; 
        'd4016: dout <= { 2'd2, 8'd024, 10'd325 }; 
        'd4017: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4018: dout <= { 2'd1, 8'd012, 10'd056 }; 
        'd4019: dout <= { 2'd2, 8'd006, 10'd309 }; 
        'd4020: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4021: dout <= { 2'd1, 8'd017, 10'd334 }; 
        'd4022: dout <= { 2'd2, 8'd018, 10'd134 }; 
        'd4023: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4024: dout <= { 2'd1, 8'd004, 10'd132 }; 
        'd4025: dout <= { 2'd2, 8'd008, 10'd011 }; 
        'd4026: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4027: dout <= { 2'd1, 8'd000, 10'd088 }; 
        'd4028: dout <= { 2'd2, 8'd017, 10'd169 }; 
        'd4029: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4030: dout <= { 2'd1, 8'd018, 10'd028 }; 
        'd4031: dout <= { 2'd2, 8'd023, 10'd115 }; 
        'd4032: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4033: dout <= { 2'd1, 8'd002, 10'd186 }; 
        'd4034: dout <= { 2'd2, 8'd013, 10'd189 }; 
        'd4035: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4036: dout <= { 2'd1, 8'd013, 10'd317 }; 
        'd4037: dout <= { 2'd2, 8'd016, 10'd030 }; 
        'd4038: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4039: dout <= { 2'd1, 8'd027, 10'd136 }; 
        'd4040: dout <= { 2'd2, 8'd029, 10'd051 }; 
        'd4041: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4042: dout <= { 2'd1, 8'd006, 10'd150 }; 
        'd4043: dout <= { 2'd2, 8'd011, 10'd116 }; 
        'd4044: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4045: dout <= { 2'd1, 8'd001, 10'd273 }; 
        'd4046: dout <= { 2'd2, 8'd012, 10'd139 }; 
        'd4047: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4048: dout <= { 2'd1, 8'd022, 10'd339 }; 
        'd4049: dout <= { 2'd2, 8'd007, 10'd205 }; 
        'd4050: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4051: dout <= { 2'd1, 8'd028, 10'd188 }; 
        'd4052: dout <= { 2'd2, 8'd005, 10'd110 }; 
        'd4053: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4054: dout <= { 2'd1, 8'd029, 10'd114 }; 
        'd4055: dout <= { 2'd2, 8'd010, 10'd051 }; 
        'd4056: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd4057: dout <= { 2'd1, 8'd026, 10'd158 }; 
        'd4058: dout <= { 2'd2, 8'd027, 10'd089 }; 
        'd4059: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd4060: dout <= { 2'd1, 8'd019, 10'd135 }; 
        'd4061: dout <= { 2'd2, 8'd015, 10'd222 }; 
        'd4062: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd4063: dout <= { 2'd1, 8'd007, 10'd037 }; 
        'd4064: dout <= { 2'd2, 8'd026, 10'd033 }; 
        'd4065: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd4066: dout <= { 2'd1, 8'd009, 10'd187 }; 
        'd4067: dout <= { 2'd2, 8'd025, 10'd102 }; 
        'd4068: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd4069: dout <= { 2'd1, 8'd023, 10'd282 }; 
        'd4070: dout <= { 2'd2, 8'd000, 10'd280 }; 
        'd4071: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd4072: dout <= { 2'd1, 8'd005, 10'd275 }; 
        'd4073: dout <= { 2'd2, 8'd004, 10'd013 }; 
        'd4074: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd4075: dout <= { 2'd1, 8'd008, 10'd211 }; 
        'd4076: dout <= { 2'd2, 8'd002, 10'd168 }; 
        'd4077: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd4078: dout <= { 2'd1, 8'd024, 10'd205 }; 
        'd4079: dout <= { 2'd2, 8'd019, 10'd170 }; 
        'd4080: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd4081: dout <= { 2'd1, 8'd003, 10'd240 }; 
        'd4082: dout <= { 2'd2, 8'd009, 10'd066 }; 
        'd4083: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd4084: dout <= { 2'd1, 8'd011, 10'd059 }; 
        'd4085: dout <= { 2'd2, 8'd014, 10'd172 }; 
        'd4086: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4087: dout <= { 2'd1, 8'd024, 10'd048 }; 
        'd4088: dout <= { 2'd2, 8'd019, 10'd118 }; 
        'd4089: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4090: dout <= { 2'd1, 8'd016, 10'd112 }; 
        'd4091: dout <= { 2'd2, 8'd014, 10'd140 }; 
        'd4092: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4093: dout <= { 2'd1, 8'd008, 10'd241 }; 
        'd4094: dout <= { 2'd2, 8'd007, 10'd002 }; 
        'd4095: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4096: dout <= { 2'd1, 8'd005, 10'd353 }; 
        'd4097: dout <= { 2'd2, 8'd011, 10'd294 }; 
        'd4098: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4099: dout <= { 2'd1, 8'd021, 10'd040 }; 
        'd4100: dout <= { 2'd2, 8'd003, 10'd217 }; 
        'd4101: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4102: dout <= { 2'd1, 8'd020, 10'd176 }; 
        'd4103: dout <= { 2'd2, 8'd002, 10'd155 }; 
        'd4104: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4105: dout <= { 2'd1, 8'd019, 10'd047 }; 
        'd4106: dout <= { 2'd2, 8'd029, 10'd324 }; 
        'd4107: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4108: dout <= { 2'd1, 8'd018, 10'd262 }; 
        'd4109: dout <= { 2'd2, 8'd001, 10'd171 }; 
        'd4110: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4111: dout <= { 2'd1, 8'd025, 10'd147 }; 
        'd4112: dout <= { 2'd2, 8'd024, 10'd342 }; 
        'd4113: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4114: dout <= { 2'd1, 8'd001, 10'd211 }; 
        'd4115: dout <= { 2'd2, 8'd017, 10'd183 }; 
        'd4116: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4117: dout <= { 2'd1, 8'd002, 10'd222 }; 
        'd4118: dout <= { 2'd2, 8'd021, 10'd164 }; 
        'd4119: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4120: dout <= { 2'd1, 8'd014, 10'd320 }; 
        'd4121: dout <= { 2'd2, 8'd008, 10'd341 }; 
        'd4122: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4123: dout <= { 2'd1, 8'd000, 10'd280 }; 
        'd4124: dout <= { 2'd2, 8'd015, 10'd267 }; 
        'd4125: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4126: dout <= { 2'd1, 8'd006, 10'd305 }; 
        'd4127: dout <= { 2'd2, 8'd020, 10'd187 }; 
        'd4128: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4129: dout <= { 2'd1, 8'd017, 10'd235 }; 
        'd4130: dout <= { 2'd2, 8'd028, 10'd295 }; 
        'd4131: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4132: dout <= { 2'd1, 8'd027, 10'd300 }; 
        'd4133: dout <= { 2'd2, 8'd025, 10'd113 }; 
        'd4134: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4135: dout <= { 2'd1, 8'd010, 10'd056 }; 
        'd4136: dout <= { 2'd2, 8'd026, 10'd128 }; 
        'd4137: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4138: dout <= { 2'd1, 8'd004, 10'd095 }; 
        'd4139: dout <= { 2'd2, 8'd009, 10'd282 }; 
        'd4140: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4141: dout <= { 2'd1, 8'd026, 10'd206 }; 
        'd4142: dout <= { 2'd2, 8'd000, 10'd021 }; 
        'd4143: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4144: dout <= { 2'd1, 8'd003, 10'd012 }; 
        'd4145: dout <= { 2'd2, 8'd023, 10'd181 }; 
        'd4146: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd4147: dout <= { 2'd1, 8'd015, 10'd137 }; 
        'd4148: dout <= { 2'd2, 8'd018, 10'd233 }; 
        'd4149: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd4150: dout <= { 2'd1, 8'd022, 10'd053 }; 
        'd4151: dout <= { 2'd2, 8'd012, 10'd223 }; 
        'd4152: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd4153: dout <= { 2'd1, 8'd009, 10'd302 }; 
        'd4154: dout <= { 2'd2, 8'd016, 10'd307 }; 
        'd4155: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd4156: dout <= { 2'd1, 8'd007, 10'd192 }; 
        'd4157: dout <= { 2'd2, 8'd010, 10'd135 }; 
        'd4158: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd4159: dout <= { 2'd1, 8'd023, 10'd124 }; 
        'd4160: dout <= { 2'd2, 8'd027, 10'd307 }; 
        'd4161: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd4162: dout <= { 2'd1, 8'd028, 10'd233 }; 
        'd4163: dout <= { 2'd2, 8'd022, 10'd185 }; 
        'd4164: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd4165: dout <= { 2'd1, 8'd012, 10'd296 }; 
        'd4166: dout <= { 2'd2, 8'd006, 10'd151 }; 
        'd4167: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd4168: dout <= { 2'd1, 8'd013, 10'd028 }; 
        'd4169: dout <= { 2'd2, 8'd004, 10'd202 }; 
        'd4170: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd4171: dout <= { 2'd1, 8'd029, 10'd268 }; 
        'd4172: dout <= { 2'd2, 8'd013, 10'd196 }; 
        'd4173: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd4174: dout <= { 2'd1, 8'd011, 10'd068 }; 
        'd4175: dout <= { 2'd2, 8'd005, 10'd096 }; 
        'd4176: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4177: dout <= { 2'd1, 8'd011, 10'd356 }; 
        'd4178: dout <= { 2'd2, 8'd003, 10'd105 }; 
        'd4179: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4180: dout <= { 2'd1, 8'd002, 10'd120 }; 
        'd4181: dout <= { 2'd2, 8'd005, 10'd135 }; 
        'd4182: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4183: dout <= { 2'd1, 8'd028, 10'd010 }; 
        'd4184: dout <= { 2'd2, 8'd007, 10'd057 }; 
        'd4185: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4186: dout <= { 2'd1, 8'd029, 10'd073 }; 
        'd4187: dout <= { 2'd2, 8'd029, 10'd309 }; 
        'd4188: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4189: dout <= { 2'd1, 8'd019, 10'd064 }; 
        'd4190: dout <= { 2'd2, 8'd008, 10'd263 }; 
        'd4191: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4192: dout <= { 2'd1, 8'd017, 10'd020 }; 
        'd4193: dout <= { 2'd2, 8'd026, 10'd006 }; 
        'd4194: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4195: dout <= { 2'd1, 8'd024, 10'd284 }; 
        'd4196: dout <= { 2'd2, 8'd024, 10'd045 }; 
        'd4197: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4198: dout <= { 2'd1, 8'd026, 10'd355 }; 
        'd4199: dout <= { 2'd2, 8'd000, 10'd108 }; 
        'd4200: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4201: dout <= { 2'd1, 8'd012, 10'd222 }; 
        'd4202: dout <= { 2'd2, 8'd009, 10'd316 }; 
        'd4203: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4204: dout <= { 2'd1, 8'd020, 10'd105 }; 
        'd4205: dout <= { 2'd2, 8'd017, 10'd248 }; 
        'd4206: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4207: dout <= { 2'd1, 8'd008, 10'd262 }; 
        'd4208: dout <= { 2'd2, 8'd001, 10'd191 }; 
        'd4209: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4210: dout <= { 2'd1, 8'd001, 10'd204 }; 
        'd4211: dout <= { 2'd2, 8'd022, 10'd357 }; 
        'd4212: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4213: dout <= { 2'd1, 8'd013, 10'd161 }; 
        'd4214: dout <= { 2'd2, 8'd012, 10'd304 }; 
        'd4215: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4216: dout <= { 2'd1, 8'd010, 10'd019 }; 
        'd4217: dout <= { 2'd2, 8'd021, 10'd319 }; 
        'd4218: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4219: dout <= { 2'd1, 8'd027, 10'd208 }; 
        'd4220: dout <= { 2'd2, 8'd020, 10'd309 }; 
        'd4221: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4222: dout <= { 2'd1, 8'd009, 10'd100 }; 
        'd4223: dout <= { 2'd2, 8'd018, 10'd075 }; 
        'd4224: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4225: dout <= { 2'd1, 8'd015, 10'd006 }; 
        'd4226: dout <= { 2'd2, 8'd019, 10'd080 }; 
        'd4227: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4228: dout <= { 2'd1, 8'd006, 10'd267 }; 
        'd4229: dout <= { 2'd2, 8'd027, 10'd051 }; 
        'd4230: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4231: dout <= { 2'd1, 8'd016, 10'd050 }; 
        'd4232: dout <= { 2'd2, 8'd015, 10'd306 }; 
        'd4233: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4234: dout <= { 2'd1, 8'd022, 10'd268 }; 
        'd4235: dout <= { 2'd2, 8'd004, 10'd302 }; 
        'd4236: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd4237: dout <= { 2'd1, 8'd025, 10'd069 }; 
        'd4238: dout <= { 2'd2, 8'd028, 10'd298 }; 
        'd4239: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd4240: dout <= { 2'd1, 8'd003, 10'd025 }; 
        'd4241: dout <= { 2'd2, 8'd006, 10'd244 }; 
        'd4242: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd4243: dout <= { 2'd1, 8'd021, 10'd209 }; 
        'd4244: dout <= { 2'd2, 8'd023, 10'd127 }; 
        'd4245: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd4246: dout <= { 2'd1, 8'd004, 10'd087 }; 
        'd4247: dout <= { 2'd2, 8'd014, 10'd261 }; 
        'd4248: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd4249: dout <= { 2'd1, 8'd023, 10'd076 }; 
        'd4250: dout <= { 2'd2, 8'd016, 10'd021 }; 
        'd4251: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd4252: dout <= { 2'd1, 8'd005, 10'd069 }; 
        'd4253: dout <= { 2'd2, 8'd011, 10'd020 }; 
        'd4254: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd4255: dout <= { 2'd1, 8'd007, 10'd156 }; 
        'd4256: dout <= { 2'd2, 8'd002, 10'd012 }; 
        'd4257: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd4258: dout <= { 2'd1, 8'd014, 10'd289 }; 
        'd4259: dout <= { 2'd2, 8'd010, 10'd331 }; 
        'd4260: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd4261: dout <= { 2'd1, 8'd000, 10'd161 }; 
        'd4262: dout <= { 2'd2, 8'd025, 10'd068 }; 
        'd4263: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd4264: dout <= { 2'd1, 8'd018, 10'd234 }; 
        'd4265: dout <= { 2'd2, 8'd013, 10'd045 }; 
        'd4266: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4267: dout <= { 2'd1, 8'd029, 10'd058 }; 
        'd4268: dout <= { 2'd2, 8'd007, 10'd261 }; 
        'd4269: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4270: dout <= { 2'd1, 8'd021, 10'd126 }; 
        'd4271: dout <= { 2'd2, 8'd009, 10'd056 }; 
        'd4272: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4273: dout <= { 2'd1, 8'd020, 10'd335 }; 
        'd4274: dout <= { 2'd2, 8'd019, 10'd078 }; 
        'd4275: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4276: dout <= { 2'd1, 8'd007, 10'd122 }; 
        'd4277: dout <= { 2'd2, 8'd018, 10'd330 }; 
        'd4278: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4279: dout <= { 2'd1, 8'd024, 10'd063 }; 
        'd4280: dout <= { 2'd2, 8'd020, 10'd230 }; 
        'd4281: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4282: dout <= { 2'd1, 8'd014, 10'd141 }; 
        'd4283: dout <= { 2'd2, 8'd029, 10'd188 }; 
        'd4284: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4285: dout <= { 2'd1, 8'd015, 10'd341 }; 
        'd4286: dout <= { 2'd2, 8'd021, 10'd260 }; 
        'd4287: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4288: dout <= { 2'd1, 8'd028, 10'd254 }; 
        'd4289: dout <= { 2'd2, 8'd014, 10'd131 }; 
        'd4290: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4291: dout <= { 2'd1, 8'd010, 10'd110 }; 
        'd4292: dout <= { 2'd2, 8'd028, 10'd182 }; 
        'd4293: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4294: dout <= { 2'd1, 8'd016, 10'd211 }; 
        'd4295: dout <= { 2'd2, 8'd006, 10'd322 }; 
        'd4296: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4297: dout <= { 2'd1, 8'd008, 10'd236 }; 
        'd4298: dout <= { 2'd2, 8'd002, 10'd204 }; 
        'd4299: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4300: dout <= { 2'd1, 8'd001, 10'd043 }; 
        'd4301: dout <= { 2'd2, 8'd027, 10'd260 }; 
        'd4302: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4303: dout <= { 2'd1, 8'd002, 10'd353 }; 
        'd4304: dout <= { 2'd2, 8'd005, 10'd298 }; 
        'd4305: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4306: dout <= { 2'd1, 8'd009, 10'd120 }; 
        'd4307: dout <= { 2'd2, 8'd010, 10'd237 }; 
        'd4308: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4309: dout <= { 2'd1, 8'd018, 10'd305 }; 
        'd4310: dout <= { 2'd2, 8'd022, 10'd303 }; 
        'd4311: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4312: dout <= { 2'd1, 8'd023, 10'd206 }; 
        'd4313: dout <= { 2'd2, 8'd012, 10'd268 }; 
        'd4314: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4315: dout <= { 2'd1, 8'd000, 10'd111 }; 
        'd4316: dout <= { 2'd2, 8'd015, 10'd096 }; 
        'd4317: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4318: dout <= { 2'd1, 8'd004, 10'd142 }; 
        'd4319: dout <= { 2'd2, 8'd003, 10'd352 }; 
        'd4320: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4321: dout <= { 2'd1, 8'd026, 10'd351 }; 
        'd4322: dout <= { 2'd2, 8'd016, 10'd216 }; 
        'd4323: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4324: dout <= { 2'd1, 8'd017, 10'd293 }; 
        'd4325: dout <= { 2'd2, 8'd025, 10'd254 }; 
        'd4326: dout <= { 2'd1, 8'd020, 10'd000 }; 
        'd4327: dout <= { 2'd1, 8'd019, 10'd066 }; 
        'd4328: dout <= { 2'd2, 8'd000, 10'd151 }; 
        'd4329: dout <= { 2'd1, 8'd021, 10'd000 }; 
        'd4330: dout <= { 2'd1, 8'd022, 10'd306 }; 
        'd4331: dout <= { 2'd2, 8'd008, 10'd227 }; 
        'd4332: dout <= { 2'd1, 8'd022, 10'd000 }; 
        'd4333: dout <= { 2'd1, 8'd013, 10'd113 }; 
        'd4334: dout <= { 2'd2, 8'd024, 10'd057 }; 
        'd4335: dout <= { 2'd1, 8'd023, 10'd000 }; 
        'd4336: dout <= { 2'd1, 8'd006, 10'd070 }; 
        'd4337: dout <= { 2'd2, 8'd023, 10'd300 }; 
        'd4338: dout <= { 2'd1, 8'd024, 10'd000 }; 
        'd4339: dout <= { 2'd1, 8'd011, 10'd229 }; 
        'd4340: dout <= { 2'd2, 8'd013, 10'd129 }; 
        'd4341: dout <= { 2'd1, 8'd025, 10'd000 }; 
        'd4342: dout <= { 2'd1, 8'd025, 10'd129 }; 
        'd4343: dout <= { 2'd2, 8'd011, 10'd072 }; 
        'd4344: dout <= { 2'd1, 8'd026, 10'd000 }; 
        'd4345: dout <= { 2'd1, 8'd012, 10'd135 }; 
        'd4346: dout <= { 2'd2, 8'd004, 10'd214 }; 
        'd4347: dout <= { 2'd1, 8'd027, 10'd000 }; 
        'd4348: dout <= { 2'd1, 8'd005, 10'd125 }; 
        'd4349: dout <= { 2'd2, 8'd026, 10'd317 }; 
        'd4350: dout <= { 2'd1, 8'd028, 10'd000 }; 
        'd4351: dout <= { 2'd1, 8'd003, 10'd156 }; 
        'd4352: dout <= { 2'd2, 8'd001, 10'd071 }; 
        'd4353: dout <= { 2'd1, 8'd029, 10'd000 }; 
        'd4354: dout <= { 2'd1, 8'd027, 10'd244 }; 
        'd4355: dout <= { 2'd3, 8'd017, 10'd267 }; 
        // Q=20, BaseAddr=4356
        'd4356: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4357: dout <= { 2'd1, 8'd015, 10'd311 }; 
        'd4358: dout <= { 2'd1, 8'd008, 10'd142 }; 
        'd4359: dout <= { 2'd2, 8'd002, 10'd161 }; 
        'd4360: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4361: dout <= { 2'd1, 8'd000, 10'd290 }; 
        'd4362: dout <= { 2'd1, 8'd012, 10'd174 }; 
        'd4363: dout <= { 2'd2, 8'd008, 10'd267 }; 
        'd4364: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4365: dout <= { 2'd1, 8'd017, 10'd137 }; 
        'd4366: dout <= { 2'd1, 8'd007, 10'd046 }; 
        'd4367: dout <= { 2'd2, 8'd010, 10'd004 }; 
        'd4368: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4369: dout <= { 2'd1, 8'd001, 10'd348 }; 
        'd4370: dout <= { 2'd1, 8'd016, 10'd225 }; 
        'd4371: dout <= { 2'd2, 8'd019, 10'd236 }; 
        'd4372: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4373: dout <= { 2'd1, 8'd012, 10'd058 }; 
        'd4374: dout <= { 2'd1, 8'd017, 10'd161 }; 
        'd4375: dout <= { 2'd2, 8'd004, 10'd313 }; 
        'd4376: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4377: dout <= { 2'd1, 8'd007, 10'd096 }; 
        'd4378: dout <= { 2'd1, 8'd005, 10'd121 }; 
        'd4379: dout <= { 2'd2, 8'd003, 10'd184 }; 
        'd4380: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4381: dout <= { 2'd1, 8'd014, 10'd185 }; 
        'd4382: dout <= { 2'd1, 8'd009, 10'd315 }; 
        'd4383: dout <= { 2'd2, 8'd015, 10'd124 }; 
        'd4384: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4385: dout <= { 2'd1, 8'd010, 10'd153 }; 
        'd4386: dout <= { 2'd1, 8'd002, 10'd317 }; 
        'd4387: dout <= { 2'd2, 8'd014, 10'd357 }; 
        'd4388: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4389: dout <= { 2'd1, 8'd008, 10'd121 }; 
        'd4390: dout <= { 2'd1, 8'd013, 10'd030 }; 
        'd4391: dout <= { 2'd2, 8'd001, 10'd188 }; 
        'd4392: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4393: dout <= { 2'd1, 8'd006, 10'd145 }; 
        'd4394: dout <= { 2'd1, 8'd004, 10'd013 }; 
        'd4395: dout <= { 2'd2, 8'd007, 10'd296 }; 
        'd4396: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4397: dout <= { 2'd1, 8'd016, 10'd085 }; 
        'd4398: dout <= { 2'd1, 8'd010, 10'd097 }; 
        'd4399: dout <= { 2'd2, 8'd013, 10'd213 }; 
        'd4400: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4401: dout <= { 2'd1, 8'd013, 10'd230 }; 
        'd4402: dout <= { 2'd1, 8'd019, 10'd308 }; 
        'd4403: dout <= { 2'd2, 8'd011, 10'd174 }; 
        'd4404: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4405: dout <= { 2'd1, 8'd005, 10'd243 }; 
        'd4406: dout <= { 2'd1, 8'd006, 10'd164 }; 
        'd4407: dout <= { 2'd2, 8'd005, 10'd300 }; 
        'd4408: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4409: dout <= { 2'd1, 8'd003, 10'd067 }; 
        'd4410: dout <= { 2'd1, 8'd003, 10'd296 }; 
        'd4411: dout <= { 2'd2, 8'd009, 10'd176 }; 
        'd4412: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4413: dout <= { 2'd1, 8'd009, 10'd229 }; 
        'd4414: dout <= { 2'd1, 8'd015, 10'd201 }; 
        'd4415: dout <= { 2'd2, 8'd012, 10'd106 }; 
        'd4416: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4417: dout <= { 2'd1, 8'd019, 10'd078 }; 
        'd4418: dout <= { 2'd1, 8'd000, 10'd196 }; 
        'd4419: dout <= { 2'd2, 8'd017, 10'd336 }; 
        'd4420: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4421: dout <= { 2'd1, 8'd004, 10'd082 }; 
        'd4422: dout <= { 2'd1, 8'd011, 10'd059 }; 
        'd4423: dout <= { 2'd2, 8'd018, 10'd299 }; 
        'd4424: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4425: dout <= { 2'd1, 8'd002, 10'd074 }; 
        'd4426: dout <= { 2'd1, 8'd001, 10'd119 }; 
        'd4427: dout <= { 2'd2, 8'd000, 10'd231 }; 
        'd4428: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4429: dout <= { 2'd1, 8'd011, 10'd339 }; 
        'd4430: dout <= { 2'd1, 8'd014, 10'd300 }; 
        'd4431: dout <= { 2'd2, 8'd016, 10'd329 }; 
        'd4432: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4433: dout <= { 2'd1, 8'd018, 10'd136 }; 
        'd4434: dout <= { 2'd1, 8'd018, 10'd295 }; 
        'd4435: dout <= { 2'd2, 8'd006, 10'd189 }; 
        'd4436: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4437: dout <= { 2'd1, 8'd016, 10'd257 }; 
        'd4438: dout <= { 2'd2, 8'd006, 10'd308 }; 
        'd4439: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4440: dout <= { 2'd1, 8'd004, 10'd075 }; 
        'd4441: dout <= { 2'd2, 8'd016, 10'd217 }; 
        'd4442: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4443: dout <= { 2'd1, 8'd010, 10'd006 }; 
        'd4444: dout <= { 2'd2, 8'd004, 10'd095 }; 
        'd4445: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4446: dout <= { 2'd1, 8'd007, 10'd301 }; 
        'd4447: dout <= { 2'd2, 8'd007, 10'd159 }; 
        'd4448: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4449: dout <= { 2'd1, 8'd018, 10'd335 }; 
        'd4450: dout <= { 2'd2, 8'd019, 10'd037 }; 
        'd4451: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4452: dout <= { 2'd1, 8'd000, 10'd312 }; 
        'd4453: dout <= { 2'd2, 8'd010, 10'd143 }; 
        'd4454: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4455: dout <= { 2'd1, 8'd003, 10'd117 }; 
        'd4456: dout <= { 2'd2, 8'd011, 10'd065 }; 
        'd4457: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4458: dout <= { 2'd1, 8'd019, 10'd051 }; 
        'd4459: dout <= { 2'd2, 8'd005, 10'd273 }; 
        'd4460: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4461: dout <= { 2'd1, 8'd017, 10'd330 }; 
        'd4462: dout <= { 2'd2, 8'd013, 10'd125 }; 
        'd4463: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4464: dout <= { 2'd1, 8'd008, 10'd079 }; 
        'd4465: dout <= { 2'd2, 8'd002, 10'd261 }; 
        'd4466: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4467: dout <= { 2'd1, 8'd001, 10'd328 }; 
        'd4468: dout <= { 2'd2, 8'd015, 10'd026 }; 
        'd4469: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4470: dout <= { 2'd1, 8'd005, 10'd238 }; 
        'd4471: dout <= { 2'd2, 8'd014, 10'd102 }; 
        'd4472: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4473: dout <= { 2'd1, 8'd006, 10'd298 }; 
        'd4474: dout <= { 2'd2, 8'd012, 10'd344 }; 
        'd4475: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4476: dout <= { 2'd1, 8'd009, 10'd098 }; 
        'd4477: dout <= { 2'd2, 8'd009, 10'd193 }; 
        'd4478: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4479: dout <= { 2'd1, 8'd011, 10'd178 }; 
        'd4480: dout <= { 2'd2, 8'd000, 10'd121 }; 
        'd4481: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4482: dout <= { 2'd1, 8'd012, 10'd231 }; 
        'd4483: dout <= { 2'd2, 8'd001, 10'd049 }; 
        'd4484: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4485: dout <= { 2'd1, 8'd015, 10'd160 }; 
        'd4486: dout <= { 2'd2, 8'd003, 10'd208 }; 
        'd4487: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4488: dout <= { 2'd1, 8'd013, 10'd048 }; 
        'd4489: dout <= { 2'd2, 8'd017, 10'd155 }; 
        'd4490: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4491: dout <= { 2'd1, 8'd002, 10'd190 }; 
        'd4492: dout <= { 2'd2, 8'd018, 10'd309 }; 
        'd4493: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4494: dout <= { 2'd1, 8'd014, 10'd189 }; 
        'd4495: dout <= { 2'd2, 8'd008, 10'd197 }; 
        'd4496: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4497: dout <= { 2'd1, 8'd016, 10'd159 }; 
        'd4498: dout <= { 2'd2, 8'd006, 10'd306 }; 
        'd4499: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4500: dout <= { 2'd1, 8'd013, 10'd028 }; 
        'd4501: dout <= { 2'd2, 8'd009, 10'd095 }; 
        'd4502: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4503: dout <= { 2'd1, 8'd010, 10'd042 }; 
        'd4504: dout <= { 2'd2, 8'd014, 10'd201 }; 
        'd4505: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4506: dout <= { 2'd1, 8'd002, 10'd281 }; 
        'd4507: dout <= { 2'd2, 8'd001, 10'd080 }; 
        'd4508: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4509: dout <= { 2'd1, 8'd005, 10'd300 }; 
        'd4510: dout <= { 2'd2, 8'd004, 10'd026 }; 
        'd4511: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4512: dout <= { 2'd1, 8'd011, 10'd262 }; 
        'd4513: dout <= { 2'd2, 8'd003, 10'd289 }; 
        'd4514: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4515: dout <= { 2'd1, 8'd012, 10'd008 }; 
        'd4516: dout <= { 2'd2, 8'd012, 10'd101 }; 
        'd4517: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4518: dout <= { 2'd1, 8'd015, 10'd093 }; 
        'd4519: dout <= { 2'd2, 8'd015, 10'd123 }; 
        'd4520: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4521: dout <= { 2'd1, 8'd017, 10'd024 }; 
        'd4522: dout <= { 2'd2, 8'd011, 10'd064 }; 
        'd4523: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4524: dout <= { 2'd1, 8'd006, 10'd128 }; 
        'd4525: dout <= { 2'd2, 8'd010, 10'd171 }; 
        'd4526: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4527: dout <= { 2'd1, 8'd009, 10'd062 }; 
        'd4528: dout <= { 2'd2, 8'd000, 10'd037 }; 
        'd4529: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4530: dout <= { 2'd1, 8'd004, 10'd147 }; 
        'd4531: dout <= { 2'd2, 8'd008, 10'd097 }; 
        'd4532: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4533: dout <= { 2'd1, 8'd008, 10'd326 }; 
        'd4534: dout <= { 2'd2, 8'd019, 10'd144 }; 
        'd4535: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4536: dout <= { 2'd1, 8'd003, 10'd112 }; 
        'd4537: dout <= { 2'd2, 8'd016, 10'd180 }; 
        'd4538: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4539: dout <= { 2'd1, 8'd007, 10'd043 }; 
        'd4540: dout <= { 2'd2, 8'd013, 10'd186 }; 
        'd4541: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4542: dout <= { 2'd1, 8'd014, 10'd068 }; 
        'd4543: dout <= { 2'd2, 8'd002, 10'd235 }; 
        'd4544: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4545: dout <= { 2'd1, 8'd018, 10'd234 }; 
        'd4546: dout <= { 2'd2, 8'd005, 10'd114 }; 
        'd4547: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4548: dout <= { 2'd1, 8'd000, 10'd238 }; 
        'd4549: dout <= { 2'd2, 8'd017, 10'd195 }; 
        'd4550: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4551: dout <= { 2'd1, 8'd019, 10'd092 }; 
        'd4552: dout <= { 2'd2, 8'd018, 10'd202 }; 
        'd4553: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4554: dout <= { 2'd1, 8'd001, 10'd307 }; 
        'd4555: dout <= { 2'd2, 8'd007, 10'd176 }; 
        'd4556: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4557: dout <= { 2'd1, 8'd008, 10'd107 }; 
        'd4558: dout <= { 2'd2, 8'd006, 10'd253 }; 
        'd4559: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4560: dout <= { 2'd1, 8'd006, 10'd065 }; 
        'd4561: dout <= { 2'd2, 8'd005, 10'd007 }; 
        'd4562: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4563: dout <= { 2'd1, 8'd019, 10'd115 }; 
        'd4564: dout <= { 2'd2, 8'd011, 10'd043 }; 
        'd4565: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4566: dout <= { 2'd1, 8'd003, 10'd173 }; 
        'd4567: dout <= { 2'd2, 8'd001, 10'd053 }; 
        'd4568: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4569: dout <= { 2'd1, 8'd014, 10'd277 }; 
        'd4570: dout <= { 2'd2, 8'd007, 10'd332 }; 
        'd4571: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4572: dout <= { 2'd1, 8'd017, 10'd291 }; 
        'd4573: dout <= { 2'd2, 8'd019, 10'd016 }; 
        'd4574: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4575: dout <= { 2'd1, 8'd001, 10'd291 }; 
        'd4576: dout <= { 2'd2, 8'd012, 10'd246 }; 
        'd4577: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4578: dout <= { 2'd1, 8'd016, 10'd317 }; 
        'd4579: dout <= { 2'd2, 8'd016, 10'd237 }; 
        'd4580: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4581: dout <= { 2'd1, 8'd010, 10'd196 }; 
        'd4582: dout <= { 2'd2, 8'd018, 10'd020 }; 
        'd4583: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4584: dout <= { 2'd1, 8'd011, 10'd010 }; 
        'd4585: dout <= { 2'd2, 8'd014, 10'd154 }; 
        'd4586: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4587: dout <= { 2'd1, 8'd007, 10'd050 }; 
        'd4588: dout <= { 2'd2, 8'd008, 10'd246 }; 
        'd4589: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4590: dout <= { 2'd1, 8'd004, 10'd179 }; 
        'd4591: dout <= { 2'd2, 8'd015, 10'd061 }; 
        'd4592: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4593: dout <= { 2'd1, 8'd002, 10'd349 }; 
        'd4594: dout <= { 2'd2, 8'd009, 10'd143 }; 
        'd4595: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4596: dout <= { 2'd1, 8'd012, 10'd080 }; 
        'd4597: dout <= { 2'd2, 8'd013, 10'd050 }; 
        'd4598: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4599: dout <= { 2'd1, 8'd013, 10'd047 }; 
        'd4600: dout <= { 2'd2, 8'd004, 10'd248 }; 
        'd4601: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4602: dout <= { 2'd1, 8'd015, 10'd227 }; 
        'd4603: dout <= { 2'd2, 8'd010, 10'd220 }; 
        'd4604: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4605: dout <= { 2'd1, 8'd005, 10'd246 }; 
        'd4606: dout <= { 2'd2, 8'd002, 10'd242 }; 
        'd4607: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4608: dout <= { 2'd1, 8'd018, 10'd288 }; 
        'd4609: dout <= { 2'd2, 8'd000, 10'd030 }; 
        'd4610: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4611: dout <= { 2'd1, 8'd009, 10'd325 }; 
        'd4612: dout <= { 2'd2, 8'd017, 10'd120 }; 
        'd4613: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4614: dout <= { 2'd1, 8'd000, 10'd063 }; 
        'd4615: dout <= { 2'd2, 8'd003, 10'd245 }; 
        'd4616: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4617: dout <= { 2'd1, 8'd009, 10'd168 }; 
        'd4618: dout <= { 2'd2, 8'd011, 10'd151 }; 
        'd4619: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4620: dout <= { 2'd1, 8'd017, 10'd177 }; 
        'd4621: dout <= { 2'd2, 8'd004, 10'd161 }; 
        'd4622: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4623: dout <= { 2'd1, 8'd008, 10'd151 }; 
        'd4624: dout <= { 2'd2, 8'd003, 10'd029 }; 
        'd4625: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4626: dout <= { 2'd1, 8'd018, 10'd162 }; 
        'd4627: dout <= { 2'd2, 8'd000, 10'd022 }; 
        'd4628: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4629: dout <= { 2'd1, 8'd006, 10'd311 }; 
        'd4630: dout <= { 2'd2, 8'd015, 10'd332 }; 
        'd4631: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4632: dout <= { 2'd1, 8'd015, 10'd244 }; 
        'd4633: dout <= { 2'd2, 8'd014, 10'd054 }; 
        'd4634: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4635: dout <= { 2'd1, 8'd001, 10'd074 }; 
        'd4636: dout <= { 2'd2, 8'd007, 10'd342 }; 
        'd4637: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4638: dout <= { 2'd1, 8'd013, 10'd221 }; 
        'd4639: dout <= { 2'd2, 8'd012, 10'd096 }; 
        'd4640: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4641: dout <= { 2'd1, 8'd007, 10'd105 }; 
        'd4642: dout <= { 2'd2, 8'd009, 10'd082 }; 
        'd4643: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4644: dout <= { 2'd1, 8'd019, 10'd105 }; 
        'd4645: dout <= { 2'd2, 8'd005, 10'd103 }; 
        'd4646: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4647: dout <= { 2'd1, 8'd003, 10'd200 }; 
        'd4648: dout <= { 2'd2, 8'd008, 10'd319 }; 
        'd4649: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4650: dout <= { 2'd1, 8'd000, 10'd336 }; 
        'd4651: dout <= { 2'd2, 8'd002, 10'd181 }; 
        'd4652: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4653: dout <= { 2'd1, 8'd014, 10'd184 }; 
        'd4654: dout <= { 2'd2, 8'd001, 10'd226 }; 
        'd4655: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4656: dout <= { 2'd1, 8'd004, 10'd058 }; 
        'd4657: dout <= { 2'd2, 8'd010, 10'd352 }; 
        'd4658: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4659: dout <= { 2'd1, 8'd005, 10'd098 }; 
        'd4660: dout <= { 2'd2, 8'd013, 10'd180 }; 
        'd4661: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4662: dout <= { 2'd1, 8'd011, 10'd216 }; 
        'd4663: dout <= { 2'd2, 8'd006, 10'd003 }; 
        'd4664: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4665: dout <= { 2'd1, 8'd010, 10'd148 }; 
        'd4666: dout <= { 2'd2, 8'd016, 10'd089 }; 
        'd4667: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4668: dout <= { 2'd1, 8'd012, 10'd232 }; 
        'd4669: dout <= { 2'd2, 8'd018, 10'd160 }; 
        'd4670: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4671: dout <= { 2'd1, 8'd002, 10'd088 }; 
        'd4672: dout <= { 2'd2, 8'd017, 10'd238 }; 
        'd4673: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4674: dout <= { 2'd1, 8'd016, 10'd286 }; 
        'd4675: dout <= { 2'd2, 8'd019, 10'd069 }; 
        'd4676: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4677: dout <= { 2'd1, 8'd010, 10'd048 }; 
        'd4678: dout <= { 2'd2, 8'd012, 10'd128 }; 
        'd4679: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4680: dout <= { 2'd1, 8'd002, 10'd103 }; 
        'd4681: dout <= { 2'd2, 8'd019, 10'd329 }; 
        'd4682: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4683: dout <= { 2'd1, 8'd017, 10'd229 }; 
        'd4684: dout <= { 2'd2, 8'd010, 10'd243 }; 
        'd4685: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4686: dout <= { 2'd1, 8'd008, 10'd061 }; 
        'd4687: dout <= { 2'd2, 8'd013, 10'd345 }; 
        'd4688: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4689: dout <= { 2'd1, 8'd019, 10'd207 }; 
        'd4690: dout <= { 2'd2, 8'd017, 10'd051 }; 
        'd4691: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4692: dout <= { 2'd1, 8'd016, 10'd145 }; 
        'd4693: dout <= { 2'd2, 8'd002, 10'd118 }; 
        'd4694: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4695: dout <= { 2'd1, 8'd015, 10'd019 }; 
        'd4696: dout <= { 2'd2, 8'd006, 10'd061 }; 
        'd4697: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4698: dout <= { 2'd1, 8'd011, 10'd345 }; 
        'd4699: dout <= { 2'd2, 8'd008, 10'd227 }; 
        'd4700: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4701: dout <= { 2'd1, 8'd018, 10'd230 }; 
        'd4702: dout <= { 2'd2, 8'd001, 10'd112 }; 
        'd4703: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4704: dout <= { 2'd1, 8'd000, 10'd206 }; 
        'd4705: dout <= { 2'd2, 8'd000, 10'd214 }; 
        'd4706: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4707: dout <= { 2'd1, 8'd005, 10'd291 }; 
        'd4708: dout <= { 2'd2, 8'd014, 10'd023 }; 
        'd4709: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4710: dout <= { 2'd1, 8'd014, 10'd107 }; 
        'd4711: dout <= { 2'd2, 8'd018, 10'd277 }; 
        'd4712: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4713: dout <= { 2'd1, 8'd013, 10'd189 }; 
        'd4714: dout <= { 2'd2, 8'd011, 10'd273 }; 
        'd4715: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4716: dout <= { 2'd1, 8'd007, 10'd285 }; 
        'd4717: dout <= { 2'd2, 8'd015, 10'd079 }; 
        'd4718: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4719: dout <= { 2'd1, 8'd003, 10'd070 }; 
        'd4720: dout <= { 2'd2, 8'd005, 10'd016 }; 
        'd4721: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4722: dout <= { 2'd1, 8'd001, 10'd330 }; 
        'd4723: dout <= { 2'd2, 8'd003, 10'd259 }; 
        'd4724: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4725: dout <= { 2'd1, 8'd009, 10'd318 }; 
        'd4726: dout <= { 2'd2, 8'd009, 10'd228 }; 
        'd4727: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4728: dout <= { 2'd1, 8'd006, 10'd242 }; 
        'd4729: dout <= { 2'd2, 8'd016, 10'd044 }; 
        'd4730: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4731: dout <= { 2'd1, 8'd012, 10'd354 }; 
        'd4732: dout <= { 2'd2, 8'd004, 10'd309 }; 
        'd4733: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4734: dout <= { 2'd1, 8'd004, 10'd338 }; 
        'd4735: dout <= { 2'd2, 8'd007, 10'd356 }; 
        'd4736: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4737: dout <= { 2'd1, 8'd018, 10'd317 }; 
        'd4738: dout <= { 2'd2, 8'd011, 10'd097 }; 
        'd4739: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4740: dout <= { 2'd1, 8'd017, 10'd155 }; 
        'd4741: dout <= { 2'd2, 8'd000, 10'd348 }; 
        'd4742: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4743: dout <= { 2'd1, 8'd010, 10'd135 }; 
        'd4744: dout <= { 2'd2, 8'd002, 10'd353 }; 
        'd4745: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4746: dout <= { 2'd1, 8'd013, 10'd056 }; 
        'd4747: dout <= { 2'd2, 8'd004, 10'd180 }; 
        'd4748: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4749: dout <= { 2'd1, 8'd014, 10'd184 }; 
        'd4750: dout <= { 2'd2, 8'd017, 10'd032 }; 
        'd4751: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4752: dout <= { 2'd1, 8'd015, 10'd067 }; 
        'd4753: dout <= { 2'd2, 8'd010, 10'd005 }; 
        'd4754: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4755: dout <= { 2'd1, 8'd009, 10'd166 }; 
        'd4756: dout <= { 2'd2, 8'd016, 10'd336 }; 
        'd4757: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4758: dout <= { 2'd1, 8'd005, 10'd125 }; 
        'd4759: dout <= { 2'd2, 8'd007, 10'd170 }; 
        'd4760: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4761: dout <= { 2'd1, 8'd002, 10'd123 }; 
        'd4762: dout <= { 2'd2, 8'd006, 10'd240 }; 
        'd4763: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4764: dout <= { 2'd1, 8'd016, 10'd210 }; 
        'd4765: dout <= { 2'd2, 8'd014, 10'd010 }; 
        'd4766: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4767: dout <= { 2'd1, 8'd008, 10'd267 }; 
        'd4768: dout <= { 2'd2, 8'd019, 10'd280 }; 
        'd4769: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4770: dout <= { 2'd1, 8'd007, 10'd331 }; 
        'd4771: dout <= { 2'd2, 8'd003, 10'd312 }; 
        'd4772: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4773: dout <= { 2'd1, 8'd004, 10'd132 }; 
        'd4774: dout <= { 2'd2, 8'd013, 10'd253 }; 
        'd4775: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4776: dout <= { 2'd1, 8'd012, 10'd210 }; 
        'd4777: dout <= { 2'd2, 8'd008, 10'd254 }; 
        'd4778: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4779: dout <= { 2'd1, 8'd003, 10'd173 }; 
        'd4780: dout <= { 2'd2, 8'd009, 10'd194 }; 
        'd4781: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4782: dout <= { 2'd1, 8'd006, 10'd265 }; 
        'd4783: dout <= { 2'd2, 8'd018, 10'd023 }; 
        'd4784: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4785: dout <= { 2'd1, 8'd000, 10'd216 }; 
        'd4786: dout <= { 2'd2, 8'd001, 10'd306 }; 
        'd4787: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4788: dout <= { 2'd1, 8'd001, 10'd198 }; 
        'd4789: dout <= { 2'd2, 8'd005, 10'd056 }; 
        'd4790: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4791: dout <= { 2'd1, 8'd019, 10'd284 }; 
        'd4792: dout <= { 2'd2, 8'd015, 10'd059 }; 
        'd4793: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4794: dout <= { 2'd1, 8'd011, 10'd325 }; 
        'd4795: dout <= { 2'd2, 8'd012, 10'd039 }; 
        'd4796: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4797: dout <= { 2'd1, 8'd014, 10'd196 }; 
        'd4798: dout <= { 2'd2, 8'd018, 10'd138 }; 
        'd4799: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4800: dout <= { 2'd1, 8'd018, 10'd161 }; 
        'd4801: dout <= { 2'd2, 8'd007, 10'd329 }; 
        'd4802: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4803: dout <= { 2'd1, 8'd011, 10'd055 }; 
        'd4804: dout <= { 2'd2, 8'd016, 10'd329 }; 
        'd4805: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4806: dout <= { 2'd1, 8'd017, 10'd072 }; 
        'd4807: dout <= { 2'd2, 8'd006, 10'd311 }; 
        'd4808: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4809: dout <= { 2'd1, 8'd006, 10'd072 }; 
        'd4810: dout <= { 2'd2, 8'd005, 10'd194 }; 
        'd4811: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4812: dout <= { 2'd1, 8'd007, 10'd195 }; 
        'd4813: dout <= { 2'd2, 8'd003, 10'd202 }; 
        'd4814: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4815: dout <= { 2'd1, 8'd019, 10'd341 }; 
        'd4816: dout <= { 2'd2, 8'd013, 10'd143 }; 
        'd4817: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4818: dout <= { 2'd1, 8'd013, 10'd086 }; 
        'd4819: dout <= { 2'd2, 8'd015, 10'd280 }; 
        'd4820: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4821: dout <= { 2'd1, 8'd002, 10'd260 }; 
        'd4822: dout <= { 2'd2, 8'd009, 10'd213 }; 
        'd4823: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4824: dout <= { 2'd1, 8'd004, 10'd151 }; 
        'd4825: dout <= { 2'd2, 8'd002, 10'd236 }; 
        'd4826: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4827: dout <= { 2'd1, 8'd005, 10'd272 }; 
        'd4828: dout <= { 2'd2, 8'd012, 10'd318 }; 
        'd4829: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4830: dout <= { 2'd1, 8'd010, 10'd018 }; 
        'd4831: dout <= { 2'd2, 8'd008, 10'd091 }; 
        'd4832: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4833: dout <= { 2'd1, 8'd015, 10'd234 }; 
        'd4834: dout <= { 2'd2, 8'd000, 10'd080 }; 
        'd4835: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4836: dout <= { 2'd1, 8'd000, 10'd034 }; 
        'd4837: dout <= { 2'd2, 8'd014, 10'd103 }; 
        'd4838: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4839: dout <= { 2'd1, 8'd001, 10'd090 }; 
        'd4840: dout <= { 2'd2, 8'd010, 10'd334 }; 
        'd4841: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4842: dout <= { 2'd1, 8'd009, 10'd133 }; 
        'd4843: dout <= { 2'd2, 8'd017, 10'd068 }; 
        'd4844: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4845: dout <= { 2'd1, 8'd003, 10'd123 }; 
        'd4846: dout <= { 2'd2, 8'd001, 10'd084 }; 
        'd4847: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4848: dout <= { 2'd1, 8'd012, 10'd298 }; 
        'd4849: dout <= { 2'd2, 8'd011, 10'd258 }; 
        'd4850: dout <= { 2'd1, 8'd018, 10'd000 }; 
        'd4851: dout <= { 2'd1, 8'd008, 10'd286 }; 
        'd4852: dout <= { 2'd2, 8'd004, 10'd214 }; 
        'd4853: dout <= { 2'd1, 8'd019, 10'd000 }; 
        'd4854: dout <= { 2'd1, 8'd016, 10'd084 }; 
        'd4855: dout <= { 2'd3, 8'd019, 10'd072 }; 
        // Q=18, BaseAddr=4856
        'd4856: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4857: dout <= { 2'd1, 8'd013, 10'd311 }; 
        'd4858: dout <= { 2'd1, 8'd007, 10'd142 }; 
        'd4859: dout <= { 2'd2, 8'd002, 10'd161 }; 
        'd4860: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4861: dout <= { 2'd1, 8'd000, 10'd290 }; 
        'd4862: dout <= { 2'd1, 8'd011, 10'd174 }; 
        'd4863: dout <= { 2'd2, 8'd007, 10'd267 }; 
        'd4864: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4865: dout <= { 2'd1, 8'd015, 10'd137 }; 
        'd4866: dout <= { 2'd1, 8'd006, 10'd046 }; 
        'd4867: dout <= { 2'd2, 8'd009, 10'd004 }; 
        'd4868: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4869: dout <= { 2'd1, 8'd001, 10'd348 }; 
        'd4870: dout <= { 2'd1, 8'd014, 10'd225 }; 
        'd4871: dout <= { 2'd2, 8'd017, 10'd236 }; 
        'd4872: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4873: dout <= { 2'd1, 8'd011, 10'd058 }; 
        'd4874: dout <= { 2'd1, 8'd016, 10'd161 }; 
        'd4875: dout <= { 2'd2, 8'd004, 10'd313 }; 
        'd4876: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4877: dout <= { 2'd1, 8'd006, 10'd096 }; 
        'd4878: dout <= { 2'd1, 8'd004, 10'd121 }; 
        'd4879: dout <= { 2'd2, 8'd003, 10'd184 }; 
        'd4880: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4881: dout <= { 2'd1, 8'd012, 10'd185 }; 
        'd4882: dout <= { 2'd1, 8'd008, 10'd315 }; 
        'd4883: dout <= { 2'd2, 8'd014, 10'd124 }; 
        'd4884: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4885: dout <= { 2'd1, 8'd007, 10'd121 }; 
        'd4886: dout <= { 2'd1, 8'd012, 10'd030 }; 
        'd4887: dout <= { 2'd2, 8'd001, 10'd188 }; 
        'd4888: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4889: dout <= { 2'd1, 8'd005, 10'd145 }; 
        'd4890: dout <= { 2'd1, 8'd002, 10'd013 }; 
        'd4891: dout <= { 2'd2, 8'd006, 10'd296 }; 
        'd4892: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4893: dout <= { 2'd1, 8'd016, 10'd085 }; 
        'd4894: dout <= { 2'd1, 8'd009, 10'd097 }; 
        'd4895: dout <= { 2'd2, 8'd012, 10'd213 }; 
        'd4896: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4897: dout <= { 2'd1, 8'd014, 10'd230 }; 
        'd4898: dout <= { 2'd1, 8'd017, 10'd308 }; 
        'd4899: dout <= { 2'd2, 8'd010, 10'd174 }; 
        'd4900: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4901: dout <= { 2'd1, 8'd008, 10'd243 }; 
        'd4902: dout <= { 2'd1, 8'd005, 10'd164 }; 
        'd4903: dout <= { 2'd2, 8'd000, 10'd300 }; 
        'd4904: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4905: dout <= { 2'd1, 8'd003, 10'd067 }; 
        'd4906: dout <= { 2'd1, 8'd001, 10'd296 }; 
        'd4907: dout <= { 2'd2, 8'd011, 10'd176 }; 
        'd4908: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4909: dout <= { 2'd1, 8'd017, 10'd078 }; 
        'd4910: dout <= { 2'd1, 8'd000, 10'd196 }; 
        'd4911: dout <= { 2'd2, 8'd015, 10'd336 }; 
        'd4912: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4913: dout <= { 2'd1, 8'd004, 10'd082 }; 
        'd4914: dout <= { 2'd1, 8'd010, 10'd059 }; 
        'd4915: dout <= { 2'd2, 8'd016, 10'd299 }; 
        'd4916: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4917: dout <= { 2'd1, 8'd009, 10'd213 }; 
        'd4918: dout <= { 2'd1, 8'd013, 10'd098 }; 
        'd4919: dout <= { 2'd2, 8'd013, 10'd242 }; 
        'd4920: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4921: dout <= { 2'd1, 8'd002, 10'd074 }; 
        'd4922: dout <= { 2'd1, 8'd003, 10'd119 }; 
        'd4923: dout <= { 2'd2, 8'd005, 10'd231 }; 
        'd4924: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4925: dout <= { 2'd1, 8'd010, 10'd131 }; 
        'd4926: dout <= { 2'd1, 8'd015, 10'd280 }; 
        'd4927: dout <= { 2'd2, 8'd008, 10'd014 }; 
        'd4928: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4929: dout <= { 2'd1, 8'd016, 10'd339 }; 
        'd4930: dout <= { 2'd2, 8'd005, 10'd300 }; 
        'd4931: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4932: dout <= { 2'd1, 8'd006, 10'd166 }; 
        'd4933: dout <= { 2'd2, 8'd014, 10'd242 }; 
        'd4934: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4935: dout <= { 2'd1, 8'd003, 10'd189 }; 
        'd4936: dout <= { 2'd2, 8'd013, 10'd092 }; 
        'd4937: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4938: dout <= { 2'd1, 8'd014, 10'd257 }; 
        'd4939: dout <= { 2'd2, 8'd006, 10'd308 }; 
        'd4940: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4941: dout <= { 2'd1, 8'd004, 10'd075 }; 
        'd4942: dout <= { 2'd2, 8'd015, 10'd217 }; 
        'd4943: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4944: dout <= { 2'd1, 8'd009, 10'd006 }; 
        'd4945: dout <= { 2'd2, 8'd003, 10'd095 }; 
        'd4946: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd4947: dout <= { 2'd1, 8'd007, 10'd301 }; 
        'd4948: dout <= { 2'd2, 8'd004, 10'd159 }; 
        'd4949: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd4950: dout <= { 2'd1, 8'd017, 10'd335 }; 
        'd4951: dout <= { 2'd2, 8'd017, 10'd037 }; 
        'd4952: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd4953: dout <= { 2'd1, 8'd000, 10'd312 }; 
        'd4954: dout <= { 2'd2, 8'd008, 10'd143 }; 
        'd4955: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd4956: dout <= { 2'd1, 8'd002, 10'd117 }; 
        'd4957: dout <= { 2'd2, 8'd009, 10'd065 }; 
        'd4958: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd4959: dout <= { 2'd1, 8'd015, 10'd051 }; 
        'd4960: dout <= { 2'd2, 8'd007, 10'd273 }; 
        'd4961: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd4962: dout <= { 2'd1, 8'd013, 10'd330 }; 
        'd4963: dout <= { 2'd2, 8'd011, 10'd125 }; 
        'd4964: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd4965: dout <= { 2'd1, 8'd008, 10'd079 }; 
        'd4966: dout <= { 2'd2, 8'd001, 10'd261 }; 
        'd4967: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd4968: dout <= { 2'd1, 8'd001, 10'd328 }; 
        'd4969: dout <= { 2'd2, 8'd012, 10'd026 }; 
        'd4970: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd4971: dout <= { 2'd1, 8'd005, 10'd238 }; 
        'd4972: dout <= { 2'd2, 8'd010, 10'd102 }; 
        'd4973: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd4974: dout <= { 2'd1, 8'd010, 10'd298 }; 
        'd4975: dout <= { 2'd2, 8'd016, 10'd344 }; 
        'd4976: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd4977: dout <= { 2'd1, 8'd011, 10'd098 }; 
        'd4978: dout <= { 2'd2, 8'd002, 10'd193 }; 
        'd4979: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd4980: dout <= { 2'd1, 8'd012, 10'd178 }; 
        'd4981: dout <= { 2'd2, 8'd000, 10'd121 }; 
        'd4982: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd4983: dout <= { 2'd1, 8'd007, 10'd231 }; 
        'd4984: dout <= { 2'd2, 8'd002, 10'd049 }; 
        'd4985: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd4986: dout <= { 2'd1, 8'd016, 10'd160 }; 
        'd4987: dout <= { 2'd2, 8'd000, 10'd208 }; 
        'd4988: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd4989: dout <= { 2'd1, 8'd010, 10'd048 }; 
        'd4990: dout <= { 2'd2, 8'd011, 10'd155 }; 
        'd4991: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd4992: dout <= { 2'd1, 8'd003, 10'd190 }; 
        'd4993: dout <= { 2'd2, 8'd017, 10'd309 }; 
        'd4994: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd4995: dout <= { 2'd1, 8'd002, 10'd189 }; 
        'd4996: dout <= { 2'd2, 8'd006, 10'd197 }; 
        'd4997: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd4998: dout <= { 2'd1, 8'd014, 10'd159 }; 
        'd4999: dout <= { 2'd2, 8'd007, 10'd306 }; 
        'd5000: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd5001: dout <= { 2'd1, 8'd012, 10'd028 }; 
        'd5002: dout <= { 2'd2, 8'd009, 10'd095 }; 
        'd5003: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd5004: dout <= { 2'd1, 8'd009, 10'd042 }; 
        'd5005: dout <= { 2'd2, 8'd013, 10'd201 }; 
        'd5006: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd5007: dout <= { 2'd1, 8'd001, 10'd281 }; 
        'd5008: dout <= { 2'd2, 8'd001, 10'd080 }; 
        'd5009: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd5010: dout <= { 2'd1, 8'd013, 10'd312 }; 
        'd5011: dout <= { 2'd2, 8'd004, 10'd033 }; 
        'd5012: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd5013: dout <= { 2'd1, 8'd005, 10'd300 }; 
        'd5014: dout <= { 2'd2, 8'd005, 10'd026 }; 
        'd5015: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd5016: dout <= { 2'd1, 8'd008, 10'd262 }; 
        'd5017: dout <= { 2'd2, 8'd008, 10'd289 }; 
        'd5018: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd5019: dout <= { 2'd1, 8'd011, 10'd008 }; 
        'd5020: dout <= { 2'd2, 8'd014, 10'd101 }; 
        'd5021: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd5022: dout <= { 2'd1, 8'd015, 10'd093 }; 
        'd5023: dout <= { 2'd2, 8'd015, 10'd123 }; 
        'd5024: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd5025: dout <= { 2'd1, 8'd017, 10'd024 }; 
        'd5026: dout <= { 2'd2, 8'd012, 10'd064 }; 
        'd5027: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd5028: dout <= { 2'd1, 8'd004, 10'd128 }; 
        'd5029: dout <= { 2'd2, 8'd010, 10'd171 }; 
        'd5030: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd5031: dout <= { 2'd1, 8'd006, 10'd062 }; 
        'd5032: dout <= { 2'd2, 8'd003, 10'd037 }; 
        'd5033: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd5034: dout <= { 2'd1, 8'd000, 10'd126 }; 
        'd5035: dout <= { 2'd2, 8'd016, 10'd319 }; 
        'd5036: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd5037: dout <= { 2'd1, 8'd010, 10'd326 }; 
        'd5038: dout <= { 2'd2, 8'd017, 10'd144 }; 
        'd5039: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd5040: dout <= { 2'd1, 8'd008, 10'd043 }; 
        'd5041: dout <= { 2'd2, 8'd011, 10'd186 }; 
        'd5042: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd5043: dout <= { 2'd1, 8'd007, 10'd068 }; 
        'd5044: dout <= { 2'd2, 8'd001, 10'd235 }; 
        'd5045: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd5046: dout <= { 2'd1, 8'd013, 10'd234 }; 
        'd5047: dout <= { 2'd2, 8'd000, 10'd114 }; 
        'd5048: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd5049: dout <= { 2'd1, 8'd002, 10'd238 }; 
        'd5050: dout <= { 2'd2, 8'd007, 10'd195 }; 
        'd5051: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd5052: dout <= { 2'd1, 8'd005, 10'd307 }; 
        'd5053: dout <= { 2'd2, 8'd016, 10'd176 }; 
        'd5054: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd5055: dout <= { 2'd1, 8'd009, 10'd107 }; 
        'd5056: dout <= { 2'd2, 8'd006, 10'd253 }; 
        'd5057: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd5058: dout <= { 2'd1, 8'd004, 10'd065 }; 
        'd5059: dout <= { 2'd2, 8'd005, 10'd007 }; 
        'd5060: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd5061: dout <= { 2'd1, 8'd001, 10'd173 }; 
        'd5062: dout <= { 2'd2, 8'd002, 10'd053 }; 
        'd5063: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd5064: dout <= { 2'd1, 8'd015, 10'd173 }; 
        'd5065: dout <= { 2'd2, 8'd008, 10'd060 }; 
        'd5066: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd5067: dout <= { 2'd1, 8'd000, 10'd291 }; 
        'd5068: dout <= { 2'd2, 8'd012, 10'd246 }; 
        'd5069: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd5070: dout <= { 2'd1, 8'd016, 10'd317 }; 
        'd5071: dout <= { 2'd2, 8'd014, 10'd237 }; 
        'd5072: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd5073: dout <= { 2'd1, 8'd012, 10'd196 }; 
        'd5074: dout <= { 2'd2, 8'd015, 10'd020 }; 
        'd5075: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd5076: dout <= { 2'd1, 8'd011, 10'd010 }; 
        'd5077: dout <= { 2'd2, 8'd010, 10'd154 }; 
        'd5078: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd5079: dout <= { 2'd1, 8'd006, 10'd050 }; 
        'd5080: dout <= { 2'd2, 8'd004, 10'd246 }; 
        'd5081: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd5082: dout <= { 2'd1, 8'd003, 10'd179 }; 
        'd5083: dout <= { 2'd2, 8'd013, 10'd061 }; 
        'd5084: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd5085: dout <= { 2'd1, 8'd014, 10'd349 }; 
        'd5086: dout <= { 2'd2, 8'd009, 10'd143 }; 
        'd5087: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd5088: dout <= { 2'd1, 8'd017, 10'd080 }; 
        'd5089: dout <= { 2'd2, 8'd003, 10'd050 }; 
        'd5090: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd5091: dout <= { 2'd1, 8'd009, 10'd047 }; 
        'd5092: dout <= { 2'd2, 8'd011, 10'd248 }; 
        'd5093: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd5094: dout <= { 2'd1, 8'd011, 10'd227 }; 
        'd5095: dout <= { 2'd2, 8'd010, 10'd220 }; 
        'd5096: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd5097: dout <= { 2'd1, 8'd005, 10'd246 }; 
        'd5098: dout <= { 2'd2, 8'd005, 10'd242 }; 
        'd5099: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd5100: dout <= { 2'd1, 8'd014, 10'd288 }; 
        'd5101: dout <= { 2'd2, 8'd001, 10'd030 }; 
        'd5102: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd5103: dout <= { 2'd1, 8'd012, 10'd063 }; 
        'd5104: dout <= { 2'd2, 8'd016, 10'd245 }; 
        'd5105: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd5106: dout <= { 2'd1, 8'd016, 10'd177 }; 
        'd5107: dout <= { 2'd2, 8'd004, 10'd161 }; 
        'd5108: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd5109: dout <= { 2'd1, 8'd006, 10'd151 }; 
        'd5110: dout <= { 2'd2, 8'd003, 10'd029 }; 
        'd5111: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd5112: dout <= { 2'd1, 8'd003, 10'd060 }; 
        'd5113: dout <= { 2'd2, 8'd002, 10'd229 }; 
        'd5114: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd5115: dout <= { 2'd1, 8'd004, 10'd129 }; 
        'd5116: dout <= { 2'd2, 8'd009, 10'd333 }; 
        'd5117: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd5118: dout <= { 2'd1, 8'd007, 10'd311 }; 
        'd5119: dout <= { 2'd2, 8'd014, 10'd332 }; 
        'd5120: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd5121: dout <= { 2'd1, 8'd002, 10'd243 }; 
        'd5122: dout <= { 2'd2, 8'd013, 10'd087 }; 
        'd5123: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd5124: dout <= { 2'd1, 8'd015, 10'd244 }; 
        'd5125: dout <= { 2'd2, 8'd012, 10'd054 }; 
        'd5126: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd5127: dout <= { 2'd1, 8'd000, 10'd074 }; 
        'd5128: dout <= { 2'd2, 8'd007, 10'd342 }; 
        'd5129: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd5130: dout <= { 2'd1, 8'd013, 10'd297 }; 
        'd5131: dout <= { 2'd2, 8'd015, 10'd220 }; 
        'd5132: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd5133: dout <= { 2'd1, 8'd017, 10'd105 }; 
        'd5134: dout <= { 2'd2, 8'd000, 10'd103 }; 
        'd5135: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd5136: dout <= { 2'd1, 8'd001, 10'd200 }; 
        'd5137: dout <= { 2'd2, 8'd006, 10'd319 }; 
        'd5138: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd5139: dout <= { 2'd1, 8'd008, 10'd336 }; 
        'd5140: dout <= { 2'd2, 8'd008, 10'd181 }; 
        'd5141: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd5142: dout <= { 2'd1, 8'd010, 10'd184 }; 
        'd5143: dout <= { 2'd2, 8'd017, 10'd226 }; 
        'd5144: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd5145: dout <= { 2'd1, 8'd004, 10'd098 }; 
        'd5146: dout <= { 2'd2, 8'd004, 10'd180 }; 
        'd5147: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd5148: dout <= { 2'd1, 8'd007, 10'd119 }; 
        'd5149: dout <= { 2'd2, 8'd000, 10'd008 }; 
        'd5150: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd5151: dout <= { 2'd1, 8'd005, 10'd088 }; 
        'd5152: dout <= { 2'd2, 8'd007, 10'd238 }; 
        'd5153: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd5154: dout <= { 2'd1, 8'd006, 10'd286 }; 
        'd5155: dout <= { 2'd2, 8'd010, 10'd069 }; 
        'd5156: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd5157: dout <= { 2'd1, 8'd001, 10'd103 }; 
        'd5158: dout <= { 2'd2, 8'd017, 10'd329 }; 
        'd5159: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd5160: dout <= { 2'd1, 8'd014, 10'd267 }; 
        'd5161: dout <= { 2'd2, 8'd006, 10'd150 }; 
        'd5162: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd5163: dout <= { 2'd1, 8'd017, 10'd081 }; 
        'd5164: dout <= { 2'd2, 8'd012, 10'd186 }; 
        'd5165: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd5166: dout <= { 2'd1, 8'd000, 10'd237 }; 
        'd5167: dout <= { 2'd2, 8'd009, 10'd038 }; 
        'd5168: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd5169: dout <= { 2'd1, 8'd016, 10'd230 }; 
        'd5170: dout <= { 2'd2, 8'd002, 10'd112 }; 
        'd5171: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd5172: dout <= { 2'd1, 8'd015, 10'd116 }; 
        'd5173: dout <= { 2'd2, 8'd014, 10'd041 }; 
        'd5174: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd5175: dout <= { 2'd1, 8'd002, 10'd206 }; 
        'd5176: dout <= { 2'd2, 8'd001, 10'd214 }; 
        'd5177: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd5178: dout <= { 2'd1, 8'd011, 10'd284 }; 
        'd5179: dout <= { 2'd2, 8'd013, 10'd051 }; 
        'd5180: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd5181: dout <= { 2'd1, 8'd008, 10'd341 }; 
        'd5182: dout <= { 2'd2, 8'd011, 10'd184 }; 
        'd5183: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd5184: dout <= { 2'd1, 8'd013, 10'd107 }; 
        'd5185: dout <= { 2'd2, 8'd016, 10'd277 }; 
        'd5186: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd5187: dout <= { 2'd1, 8'd010, 10'd285 }; 
        'd5188: dout <= { 2'd2, 8'd015, 10'd079 }; 
        'd5189: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd5190: dout <= { 2'd1, 8'd003, 10'd070 }; 
        'd5191: dout <= { 2'd2, 8'd005, 10'd016 }; 
        'd5192: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd5193: dout <= { 2'd1, 8'd009, 10'd330 }; 
        'd5194: dout <= { 2'd2, 8'd003, 10'd259 }; 
        'd5195: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd5196: dout <= { 2'd1, 8'd012, 10'd252 }; 
        'd5197: dout <= { 2'd2, 8'd008, 10'd354 }; 
        'd5198: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd5199: dout <= { 2'd1, 8'd003, 10'd176 }; 
        'd5200: dout <= { 2'd2, 8'd010, 10'd260 }; 
        'd5201: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd5202: dout <= { 2'd1, 8'd002, 10'd289 }; 
        'd5203: dout <= { 2'd2, 8'd008, 10'd117 }; 
        'd5204: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd5205: dout <= { 2'd1, 8'd012, 10'd354 }; 
        'd5206: dout <= { 2'd2, 8'd003, 10'd309 }; 
        'd5207: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd5208: dout <= { 2'd1, 8'd016, 10'd317 }; 
        'd5209: dout <= { 2'd2, 8'd011, 10'd097 }; 
        'd5210: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd5211: dout <= { 2'd1, 8'd015, 10'd155 }; 
        'd5212: dout <= { 2'd2, 8'd000, 10'd348 }; 
        'd5213: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd5214: dout <= { 2'd1, 8'd014, 10'd066 }; 
        'd5215: dout <= { 2'd2, 8'd006, 10'd145 }; 
        'd5216: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd5217: dout <= { 2'd1, 8'd010, 10'd056 }; 
        'd5218: dout <= { 2'd2, 8'd004, 10'd180 }; 
        'd5219: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd5220: dout <= { 2'd1, 8'd004, 10'd223 }; 
        'd5221: dout <= { 2'd2, 8'd015, 10'd293 }; 
        'd5222: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd5223: dout <= { 2'd1, 8'd007, 10'd125 }; 
        'd5224: dout <= { 2'd2, 8'd007, 10'd170 }; 
        'd5225: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd5226: dout <= { 2'd1, 8'd017, 10'd137 }; 
        'd5227: dout <= { 2'd2, 8'd013, 10'd170 }; 
        'd5228: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd5229: dout <= { 2'd1, 8'd008, 10'd066 }; 
        'd5230: dout <= { 2'd2, 8'd001, 10'd296 }; 
        'd5231: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd5232: dout <= { 2'd1, 8'd001, 10'd036 }; 
        'd5233: dout <= { 2'd2, 8'd012, 10'd217 }; 
        'd5234: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd5235: dout <= { 2'd1, 8'd011, 10'd210 }; 
        'd5236: dout <= { 2'd2, 8'd009, 10'd254 }; 
        'd5237: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd5238: dout <= { 2'd1, 8'd006, 10'd279 }; 
        'd5239: dout <= { 2'd2, 8'd005, 10'd211 }; 
        'd5240: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd5241: dout <= { 2'd1, 8'd005, 10'd173 }; 
        'd5242: dout <= { 2'd2, 8'd014, 10'd194 }; 
        'd5243: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd5244: dout <= { 2'd1, 8'd009, 10'd265 }; 
        'd5245: dout <= { 2'd2, 8'd017, 10'd023 }; 
        'd5246: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd5247: dout <= { 2'd1, 8'd000, 10'd216 }; 
        'd5248: dout <= { 2'd2, 8'd002, 10'd306 }; 
        'd5249: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd5250: dout <= { 2'd1, 8'd013, 10'd243 }; 
        'd5251: dout <= { 2'd2, 8'd016, 10'd226 }; 
        'd5252: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd5253: dout <= { 2'd1, 8'd004, 10'd324 }; 
        'd5254: dout <= { 2'd2, 8'd000, 10'd094 }; 
        'd5255: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd5256: dout <= { 2'd1, 8'd014, 10'd284 }; 
        'd5257: dout <= { 2'd2, 8'd016, 10'd059 }; 
        'd5258: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd5259: dout <= { 2'd1, 8'd015, 10'd317 }; 
        'd5260: dout <= { 2'd2, 8'd009, 10'd342 }; 
        'd5261: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd5262: dout <= { 2'd1, 8'd012, 10'd196 }; 
        'd5263: dout <= { 2'd2, 8'd015, 10'd138 }; 
        'd5264: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd5265: dout <= { 2'd1, 8'd011, 10'd123 }; 
        'd5266: dout <= { 2'd2, 8'd012, 10'd352 }; 
        'd5267: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd5268: dout <= { 2'd1, 8'd000, 10'd058 }; 
        'd5269: dout <= { 2'd2, 8'd008, 10'd082 }; 
        'd5270: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd5271: dout <= { 2'd1, 8'd005, 10'd351 }; 
        'd5272: dout <= { 2'd2, 8'd010, 10'd224 }; 
        'd5273: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd5274: dout <= { 2'd1, 8'd017, 10'd072 }; 
        'd5275: dout <= { 2'd2, 8'd005, 10'd311 }; 
        'd5276: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd5277: dout <= { 2'd1, 8'd007, 10'd072 }; 
        'd5278: dout <= { 2'd2, 8'd004, 10'd194 }; 
        'd5279: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd5280: dout <= { 2'd1, 8'd006, 10'd195 }; 
        'd5281: dout <= { 2'd2, 8'd003, 10'd202 }; 
        'd5282: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd5283: dout <= { 2'd1, 8'd013, 10'd286 }; 
        'd5284: dout <= { 2'd2, 8'd007, 10'd127 }; 
        'd5285: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd5286: dout <= { 2'd1, 8'd002, 10'd260 }; 
        'd5287: dout <= { 2'd2, 8'd011, 10'd213 }; 
        'd5288: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd5289: dout <= { 2'd1, 8'd003, 10'd169 }; 
        'd5290: dout <= { 2'd2, 8'd013, 10'd035 }; 
        'd5291: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd5292: dout <= { 2'd1, 8'd010, 10'd156 }; 
        'd5293: dout <= { 2'd2, 8'd006, 10'd145 }; 
        'd5294: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd5295: dout <= { 2'd1, 8'd009, 10'd181 }; 
        'd5296: dout <= { 2'd2, 8'd001, 10'd036 }; 
        'd5297: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd5298: dout <= { 2'd1, 8'd008, 10'd346 }; 
        'd5299: dout <= { 2'd2, 8'd017, 10'd032 }; 
        'd5300: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd5301: dout <= { 2'd1, 8'd016, 10'd035 }; 
        'd5302: dout <= { 2'd2, 8'd014, 10'd163 }; 
        'd5303: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd5304: dout <= { 2'd1, 8'd001, 10'd234 }; 
        'd5305: dout <= { 2'd2, 8'd002, 10'd080 }; 
        'd5306: dout <= { 2'd1, 8'd000, 10'd000 }; 
        'd5307: dout <= { 2'd1, 8'd001, 10'd321 }; 
        'd5308: dout <= { 2'd2, 8'd012, 10'd088 }; 
        'd5309: dout <= { 2'd1, 8'd001, 10'd000 }; 
        'd5310: dout <= { 2'd1, 8'd009, 10'd133 }; 
        'd5311: dout <= { 2'd2, 8'd013, 10'd068 }; 
        'd5312: dout <= { 2'd1, 8'd002, 10'd000 }; 
        'd5313: dout <= { 2'd1, 8'd003, 10'd123 }; 
        'd5314: dout <= { 2'd2, 8'd002, 10'd084 }; 
        'd5315: dout <= { 2'd1, 8'd003, 10'd000 }; 
        'd5316: dout <= { 2'd1, 8'd011, 10'd311 }; 
        'd5317: dout <= { 2'd2, 8'd014, 10'd039 }; 
        'd5318: dout <= { 2'd1, 8'd004, 10'd000 }; 
        'd5319: dout <= { 2'd1, 8'd007, 10'd286 }; 
        'd5320: dout <= { 2'd2, 8'd006, 10'd214 }; 
        'd5321: dout <= { 2'd1, 8'd005, 10'd000 }; 
        'd5322: dout <= { 2'd1, 8'd005, 10'd084 }; 
        'd5323: dout <= { 2'd2, 8'd016, 10'd072 }; 
        'd5324: dout <= { 2'd1, 8'd006, 10'd000 }; 
        'd5325: dout <= { 2'd1, 8'd016, 10'd141 }; 
        'd5326: dout <= { 2'd2, 8'd008, 10'd175 }; 
        'd5327: dout <= { 2'd1, 8'd007, 10'd000 }; 
        'd5328: dout <= { 2'd1, 8'd006, 10'd293 }; 
        'd5329: dout <= { 2'd2, 8'd015, 10'd146 }; 
        'd5330: dout <= { 2'd1, 8'd008, 10'd000 }; 
        'd5331: dout <= { 2'd1, 8'd004, 10'd277 }; 
        'd5332: dout <= { 2'd2, 8'd003, 10'd075 }; 
        'd5333: dout <= { 2'd1, 8'd009, 10'd000 }; 
        'd5334: dout <= { 2'd1, 8'd014, 10'd313 }; 
        'd5335: dout <= { 2'd2, 8'd000, 10'd065 }; 
        'd5336: dout <= { 2'd1, 8'd010, 10'd000 }; 
        'd5337: dout <= { 2'd1, 8'd000, 10'd064 }; 
        'd5338: dout <= { 2'd2, 8'd010, 10'd242 }; 
        'd5339: dout <= { 2'd1, 8'd011, 10'd000 }; 
        'd5340: dout <= { 2'd1, 8'd015, 10'd197 }; 
        'd5341: dout <= { 2'd2, 8'd004, 10'd298 }; 
        'd5342: dout <= { 2'd1, 8'd012, 10'd000 }; 
        'd5343: dout <= { 2'd1, 8'd017, 10'd198 }; 
        'd5344: dout <= { 2'd2, 8'd007, 10'd078 }; 
        'd5345: dout <= { 2'd1, 8'd013, 10'd000 }; 
        'd5346: dout <= { 2'd1, 8'd013, 10'd313 }; 
        'd5347: dout <= { 2'd2, 8'd017, 10'd258 }; 
        'd5348: dout <= { 2'd1, 8'd014, 10'd000 }; 
        'd5349: dout <= { 2'd1, 8'd012, 10'd085 }; 
        'd5350: dout <= { 2'd2, 8'd001, 10'd300 }; 
        'd5351: dout <= { 2'd1, 8'd015, 10'd000 }; 
        'd5352: dout <= { 2'd1, 8'd002, 10'd282 }; 
        'd5353: dout <= { 2'd2, 8'd005, 10'd149 }; 
        'd5354: dout <= { 2'd1, 8'd016, 10'd000 }; 
        'd5355: dout <= { 2'd1, 8'd010, 10'd017 }; 
        'd5356: dout <= { 2'd2, 8'd009, 10'd097 }; 
        'd5357: dout <= { 2'd1, 8'd017, 10'd000 }; 
        'd5358: dout <= { 2'd1, 8'd008, 10'd188 }; 
        'd5359: dout <= { 2'd3, 8'd011, 10'd110 }; 
    endcase
end
endmodule
